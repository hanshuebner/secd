
library ieee;
use ieee.std_logic_1164.all;

package config is

  constant fep_only : std_logic := '0'; -- set to '1' to only create the FEP,
                                        -- not the SECD CPU

end;

