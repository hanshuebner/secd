
-- Automatically generated RAM initialization definitions for SECD program ../lispkit/LKIT-2/NQUEEN.LKC and argument 11


library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package secd_ram_defs is

constant RAM_SIZE : integer := 16384;
constant RAM_ADDRESS_BITS : integer := 14;
type RAM_TYPE is array (0 to (RAM_SIZE - 1)) of std_logic_vector (31 downto 0);
constant RAM_INIT : RAM_TYPE := (
 "00100000000000000000000000000000", -- 0 NIL #<SYMBOL NIL>
 "00100000000000000000000000000001", -- 1 TRUE #<SYMBOL T>
 "00100000000000000000000000000010", -- 2 FALSE #<SYMBOL F>
 "00110000000000000000000000000110", -- 3 PROG #<NUMBER 6>
 "00110000000000000000000000000010", -- 4 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 5 PROG #<SYMBOL NIL>
 "00110000000000000000000000000011", -- 6 PROG #<NUMBER 3>
 "00110000000000000000000000000001", -- 7 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 8 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 9 PROG #<NUMBER 0>
 "00000000000000100000000000001001", -- 10 PROG #<CONS 8 9>
 "00110000000000000000000000000001", -- 11 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 12 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 13 PROG #<NUMBER 1>
 "00000000000000110000000000001101", -- 14 PROG #<CONS 12 13>
 "00110000000000000000000000001110", -- 15 PROG #<NUMBER 14>
 "00110000000000000000000000001000", -- 16 PROG #<NUMBER 8>
 "00110000000000000000000000000010", -- 17 PROG #<NUMBER 2>
 "00100000000000000000000000000001", -- 18 PROG #<SYMBOL T>
 "00110000000000000000000000001001", -- 19 PROG #<NUMBER 9>
 "00000000000001001100000000000000", -- 20 PROG #<CONS 19 0>
 "00000000000001001000000000010100", -- 21 PROG #<CONS 18 20>
 "00000000000001000100000000010101", -- 22 PROG #<CONS 17 21>
 "00110000000000000000000000000001", -- 23 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 24 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 25 PROG #<NUMBER 2>
 "00000000000001100000000000011001", -- 26 PROG #<CONS 24 25>
 "00110000000000000000000000000001", -- 27 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 28 PROG #<NUMBER 0>
 "00110000000000000000000000000011", -- 29 PROG #<NUMBER 3>
 "00000000000001110000000000011101", -- 30 PROG #<CONS 28 29>
 "00110000000000000000000000001110", -- 31 PROG #<NUMBER 14>
 "00110000000000000000000000001000", -- 32 PROG #<NUMBER 8>
 "00110000000000000000000000000010", -- 33 PROG #<NUMBER 2>
 "00100000000000000000000000000001", -- 34 PROG #<SYMBOL T>
 "00110000000000000000000000001001", -- 35 PROG #<NUMBER 9>
 "00000000000010001100000000000000", -- 36 PROG #<CONS 35 0>
 "00000000000010001000000000100100", -- 37 PROG #<CONS 34 36>
 "00000000000010000100000000100101", -- 38 PROG #<CONS 33 37>
 "00110000000000000000000000000001", -- 39 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 40 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 41 PROG #<NUMBER 0>
 "00000000000010100000000000101001", -- 42 PROG #<CONS 40 41>
 "00110000000000000000000000000001", -- 43 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 44 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 45 PROG #<NUMBER 2>
 "00000000000010110000000000101101", -- 46 PROG #<CONS 44 45>
 "00110000000000000000000000001111", -- 47 PROG #<NUMBER 15>
 "00110000000000000000000000000001", -- 48 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 49 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 50 PROG #<NUMBER 1>
 "00000000000011000100000000110010", -- 51 PROG #<CONS 49 50>
 "00110000000000000000000000000001", -- 52 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 53 PROG #<NUMBER 0>
 "00110000000000000000000000000011", -- 54 PROG #<NUMBER 3>
 "00000000000011010100000000110110", -- 55 PROG #<CONS 53 54>
 "00110000000000000000000000001111", -- 56 PROG #<NUMBER 15>
 "00110000000000000000000000001110", -- 57 PROG #<NUMBER 14>
 "00110000000000000000000000001000", -- 58 PROG #<NUMBER 8>
 "00110000000000000000000000000010", -- 59 PROG #<NUMBER 2>
 "00100000000000000000000000000001", -- 60 PROG #<SYMBOL T>
 "00110000000000000000000000001001", -- 61 PROG #<NUMBER 9>
 "00000000000011110100000000000000", -- 62 PROG #<CONS 61 0>
 "00000000000011110000000000111110", -- 63 PROG #<CONS 60 62>
 "00000000000011101100000000111111", -- 64 PROG #<CONS 59 63>
 "00110000000000000000000000000001", -- 65 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 66 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 67 PROG #<NUMBER 0>
 "00000000000100001000000001000011", -- 68 PROG #<CONS 66 67>
 "00110000000000000000000000000001", -- 69 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 70 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 71 PROG #<NUMBER 2>
 "00000000000100011000000001000111", -- 72 PROG #<CONS 70 71>
 "00110000000000000000000000010000", -- 73 PROG #<NUMBER 16>
 "00110000000000000000000000000001", -- 74 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 75 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 76 PROG #<NUMBER 1>
 "00000000000100101100000001001100", -- 77 PROG #<CONS 75 76>
 "00110000000000000000000000000001", -- 78 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 79 PROG #<NUMBER 0>
 "00110000000000000000000000000011", -- 80 PROG #<NUMBER 3>
 "00000000000100111100000001010000", -- 81 PROG #<CONS 79 80>
 "00110000000000000000000000010000", -- 82 PROG #<NUMBER 16>
 "00110000000000000000000000001110", -- 83 PROG #<NUMBER 14>
 "00110000000000000000000000001000", -- 84 PROG #<NUMBER 8>
 "00110000000000000000000000000010", -- 85 PROG #<NUMBER 2>
 "00100000000000000000000000000001", -- 86 PROG #<SYMBOL T>
 "00110000000000000000000000001001", -- 87 PROG #<NUMBER 9>
 "00000000000101011100000000000000", -- 88 PROG #<CONS 87 0>
 "00000000000101011000000001011000", -- 89 PROG #<CONS 86 88>
 "00000000000101010100000001011001", -- 90 PROG #<CONS 85 89>
 "00110000000000000000000000000010", -- 91 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 92 PROG #<SYMBOL NIL>
 "00110000000000000000000000000001", -- 93 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 94 PROG #<NUMBER 0>
 "00110000000000000000000000000100", -- 95 PROG #<NUMBER 4>
 "00000000000101111000000001011111", -- 96 PROG #<CONS 94 95>
 "00110000000000000000000000001011", -- 97 PROG #<NUMBER 11>
 "00110000000000000000000000001101", -- 98 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 99 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 100 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 101 PROG #<NUMBER 2>
 "00000000000110010000000001100101", -- 102 PROG #<CONS 100 101>
 "00110000000000000000000000001101", -- 103 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 104 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 105 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 106 PROG #<NUMBER 0>
 "00000000000110100100000001101010", -- 107 PROG #<CONS 105 106>
 "00110000000000000000000000001101", -- 108 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 109 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 110 PROG #<NUMBER 1>
 "00110000000000000000000000000101", -- 111 PROG #<NUMBER 5>
 "00000000000110111000000001101111", -- 112 PROG #<CONS 110 111>
 "00110000000000000000000000000100", -- 113 PROG #<NUMBER 4>
 "00110000000000000000000000001001", -- 114 PROG #<NUMBER 9>
 "00000000000111001000000000000000", -- 115 PROG #<CONS 114 0>
 "00000000000111000100000001110011", -- 116 PROG #<CONS 113 115>
 "00000000000111000000000001110100", -- 117 PROG #<CONS 112 116>
 "00000000000110110100000001110101", -- 118 PROG #<CONS 109 117>
 "00000000000110110000000001110110", -- 119 PROG #<CONS 108 118>
 "00000000000110101100000001110111", -- 120 PROG #<CONS 107 119>
 "00000000000110100000000001111000", -- 121 PROG #<CONS 104 120>
 "00000000000110011100000001111001", -- 122 PROG #<CONS 103 121>
 "00000000000110011000000001111010", -- 123 PROG #<CONS 102 122>
 "00000000000110001100000001111011", -- 124 PROG #<CONS 99 123>
 "00000000000110001000000001111100", -- 125 PROG #<CONS 98 124>
 "00000000000110000100000001111101", -- 126 PROG #<CONS 97 125>
 "00000000000110000000000001111110", -- 127 PROG #<CONS 96 126>
 "00000000000101110100000001111111", -- 128 PROG #<CONS 93 127>
 "00000000000101110000000010000000", -- 129 PROG #<CONS 92 128>
 "00000000000101101100000010000001", -- 130 PROG #<CONS 91 129>
 "00110000000000000000000000001001", -- 131 PROG #<NUMBER 9>
 "00000000001000001100000000000000", -- 132 PROG #<CONS 131 0>
 "00000000001000001000000010000100", -- 133 PROG #<CONS 130 132>
 "00000000000101101000000010000101", -- 134 PROG #<CONS 90 133>
 "00000000000101010000000010000110", -- 135 PROG #<CONS 84 134>
 "00000000000101001100000010000111", -- 136 PROG #<CONS 83 135>
 "00000000000101001000000010001000", -- 137 PROG #<CONS 82 136>
 "00000000000101000100000010001001", -- 138 PROG #<CONS 81 137>
 "00000000000100111000000010001010", -- 139 PROG #<CONS 78 138>
 "00000000000100110100000010001011", -- 140 PROG #<CONS 77 139>
 "00000000000100101000000010001100", -- 141 PROG #<CONS 74 140>
 "00000000000100100100000010001101", -- 142 PROG #<CONS 73 141>
 "00000000000100100000000010001110", -- 143 PROG #<CONS 72 142>
 "00000000000100010100000010001111", -- 144 PROG #<CONS 69 143>
 "00000000000100010000000010010000", -- 145 PROG #<CONS 68 144>
 "00000000000100000100000010010001", -- 146 PROG #<CONS 65 145>
 "00110000000000000000000000001001", -- 147 PROG #<NUMBER 9>
 "00000000001001001100000000000000", -- 148 PROG #<CONS 147 0>
 "00000000001001001000000010010100", -- 149 PROG #<CONS 146 148>
 "00000000000100000000000010010101", -- 150 PROG #<CONS 64 149>
 "00000000000011101000000010010110", -- 151 PROG #<CONS 58 150>
 "00000000000011100100000010010111", -- 152 PROG #<CONS 57 151>
 "00000000000011100000000010011000", -- 153 PROG #<CONS 56 152>
 "00000000000011011100000010011001", -- 154 PROG #<CONS 55 153>
 "00000000000011010000000010011010", -- 155 PROG #<CONS 52 154>
 "00000000000011001100000010011011", -- 156 PROG #<CONS 51 155>
 "00000000000011000000000010011100", -- 157 PROG #<CONS 48 156>
 "00000000000010111100000010011101", -- 158 PROG #<CONS 47 157>
 "00000000000010111000000010011110", -- 159 PROG #<CONS 46 158>
 "00000000000010101100000010011111", -- 160 PROG #<CONS 43 159>
 "00000000000010101000000010100000", -- 161 PROG #<CONS 42 160>
 "00000000000010011100000010100001", -- 162 PROG #<CONS 39 161>
 "00110000000000000000000000001001", -- 163 PROG #<NUMBER 9>
 "00000000001010001100000000000000", -- 164 PROG #<CONS 163 0>
 "00000000001010001000000010100100", -- 165 PROG #<CONS 162 164>
 "00000000000010011000000010100101", -- 166 PROG #<CONS 38 165>
 "00000000000010000000000010100110", -- 167 PROG #<CONS 32 166>
 "00000000000001111100000010100111", -- 168 PROG #<CONS 31 167>
 "00000000000001111000000010101000", -- 169 PROG #<CONS 30 168>
 "00000000000001101100000010101001", -- 170 PROG #<CONS 27 169>
 "00000000000001101000000010101010", -- 171 PROG #<CONS 26 170>
 "00000000000001011100000010101011", -- 172 PROG #<CONS 23 171>
 "00110000000000000000000000000101", -- 173 PROG #<NUMBER 5>
 "00000000001010110100000000000000", -- 174 PROG #<CONS 173 0>
 "00000000001010110000000010101110", -- 175 PROG #<CONS 172 174>
 "00000000000001011000000010101111", -- 176 PROG #<CONS 22 175>
 "00000000000001000000000010110000", -- 177 PROG #<CONS 16 176>
 "00000000000000111100000010110001", -- 178 PROG #<CONS 15 177>
 "00000000000000111000000010110010", -- 179 PROG #<CONS 14 178>
 "00000000000000101100000010110011", -- 180 PROG #<CONS 11 179>
 "00000000000000101000000010110100", -- 181 PROG #<CONS 10 180>
 "00000000000000011100000010110101", -- 182 PROG #<CONS 7 181>
 "00110000000000000000000000001101", -- 183 PROG #<NUMBER 13>
 "00110000000000000000000000000011", -- 184 PROG #<NUMBER 3>
 "00110000000000000000000000000001", -- 185 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 186 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 187 PROG #<NUMBER 2>
 "00000000001011101000000010111011", -- 188 PROG #<CONS 186 187>
 "00110000000000000000000000000010", -- 189 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 190 PROG #<SYMBOL NIL>
 "00110000000000000000000000001110", -- 191 PROG #<NUMBER 14>
 "00110000000000000000000000001000", -- 192 PROG #<NUMBER 8>
 "00110000000000000000000000000010", -- 193 PROG #<NUMBER 2>
 "00100000000000000000000000000010", -- 194 PROG #<SYMBOL F>
 "00110000000000000000000000001001", -- 195 PROG #<NUMBER 9>
 "00000000001100001100000000000000", -- 196 PROG #<CONS 195 0>
 "00000000001100001000000011000100", -- 197 PROG #<CONS 194 196>
 "00000000001100000100000011000101", -- 198 PROG #<CONS 193 197>
 "00110000000000000000000000000010", -- 199 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 200 PROG #<SYMBOL NIL>
 "00110000000000000000000000000001", -- 201 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 202 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 203 PROG #<NUMBER 2>
 "00000000001100101000000011001011", -- 204 PROG #<CONS 202 203>
 "00110000000000000000000000001101", -- 205 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 206 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 207 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 208 PROG #<NUMBER 2>
 "00000000001100111100000011010000", -- 209 PROG #<CONS 207 208>
 "00110000000000000000000000001010", -- 210 PROG #<NUMBER 10>
 "00110000000000000000000000001011", -- 211 PROG #<NUMBER 11>
 "00110000000000000000000000001101", -- 212 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 213 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 214 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 215 PROG #<NUMBER 1>
 "00000000001101011000000011010111", -- 216 PROG #<CONS 214 215>
 "00110000000000000000000000001101", -- 217 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 218 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 219 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 220 PROG #<NUMBER 2>
 "00000000001101101100000011011100", -- 221 PROG #<CONS 219 220>
 "00110000000000000000000000001010", -- 222 PROG #<NUMBER 10>
 "00110000000000000000000000001010", -- 223 PROG #<NUMBER 10>
 "00110000000000000000000000001101", -- 224 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 225 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 226 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 227 PROG #<NUMBER 0>
 "00000000001110001000000011100011", -- 228 PROG #<CONS 226 227>
 "00110000000000000000000000001101", -- 229 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 230 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 231 PROG #<NUMBER 1>
 "00110000000000000000000000000110", -- 232 PROG #<NUMBER 6>
 "00000000001110011100000011101000", -- 233 PROG #<CONS 231 232>
 "00110000000000000000000000000100", -- 234 PROG #<NUMBER 4>
 "00110000000000000000000000001001", -- 235 PROG #<NUMBER 9>
 "00000000001110101100000000000000", -- 236 PROG #<CONS 235 0>
 "00000000001110101000000011101100", -- 237 PROG #<CONS 234 236>
 "00000000001110100100000011101101", -- 238 PROG #<CONS 233 237>
 "00000000001110011000000011101110", -- 239 PROG #<CONS 230 238>
 "00000000001110010100000011101111", -- 240 PROG #<CONS 229 239>
 "00000000001110010000000011110000", -- 241 PROG #<CONS 228 240>
 "00000000001110000100000011110001", -- 242 PROG #<CONS 225 241>
 "00000000001110000000000011110010", -- 243 PROG #<CONS 224 242>
 "00000000001101111100000011110011", -- 244 PROG #<CONS 223 243>
 "00000000001101111000000011110100", -- 245 PROG #<CONS 222 244>
 "00000000001101110100000011110101", -- 246 PROG #<CONS 221 245>
 "00000000001101101000000011110110", -- 247 PROG #<CONS 218 246>
 "00000000001101100100000011110111", -- 248 PROG #<CONS 217 247>
 "00000000001101100000000011111000", -- 249 PROG #<CONS 216 248>
 "00000000001101010100000011111001", -- 250 PROG #<CONS 213 249>
 "00000000001101010000000011111010", -- 251 PROG #<CONS 212 250>
 "00000000001101001100000011111011", -- 252 PROG #<CONS 211 251>
 "00000000001101001000000011111100", -- 253 PROG #<CONS 210 252>
 "00000000001101000100000011111101", -- 254 PROG #<CONS 209 253>
 "00000000001100111000000011111110", -- 255 PROG #<CONS 206 254>
 "00000000001100110100000011111111", -- 256 PROG #<CONS 205 255>
 "00000000001100110000000100000000", -- 257 PROG #<CONS 204 256>
 "00000000001100100100000100000001", -- 258 PROG #<CONS 201 257>
 "00000000001100100000000100000010", -- 259 PROG #<CONS 200 258>
 "00000000001100011100000100000011", -- 260 PROG #<CONS 199 259>
 "00110000000000000000000000000101", -- 261 PROG #<NUMBER 5>
 "00000000010000010100000000000000", -- 262 PROG #<CONS 261 0>
 "00000000010000010000000100000110", -- 263 PROG #<CONS 260 262>
 "00000000001100011000000100000111", -- 264 PROG #<CONS 198 263>
 "00000000001100000000000100001000", -- 265 PROG #<CONS 192 264>
 "00000000001011111100000100001001", -- 266 PROG #<CONS 191 265>
 "00000000001011111000000100001010", -- 267 PROG #<CONS 190 266>
 "00000000001011110100000100001011", -- 268 PROG #<CONS 189 267>
 "00000000001011110000000100001100", -- 269 PROG #<CONS 188 268>
 "00000000001011100100000100001101", -- 270 PROG #<CONS 185 269>
 "00110000000000000000000000001101", -- 271 PROG #<NUMBER 13>
 "00110000000000000000000000000011", -- 272 PROG #<NUMBER 3>
 "00110000000000000000000000000001", -- 273 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 274 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 275 PROG #<NUMBER 0>
 "00000000010001001000000100010011", -- 276 PROG #<CONS 274 275>
 "00110000000000000000000000000001", -- 277 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 278 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 279 PROG #<NUMBER 1>
 "00000000010001011000000100010111", -- 280 PROG #<CONS 278 279>
 "00110000000000000000000000001110", -- 281 PROG #<NUMBER 14>
 "00110000000000000000000000001000", -- 282 PROG #<NUMBER 8>
 "00110000000000000000000000000001", -- 283 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 284 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 285 PROG #<NUMBER 2>
 "00000000010001110000000100011101", -- 286 PROG #<CONS 284 285>
 "00110000000000000000000000001001", -- 287 PROG #<NUMBER 9>
 "00000000010001111100000000000000", -- 288 PROG #<CONS 287 0>
 "00000000010001111000000100100000", -- 289 PROG #<CONS 286 288>
 "00000000010001101100000100100001", -- 290 PROG #<CONS 283 289>
 "00110000000000000000000000000010", -- 291 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 292 PROG #<SYMBOL NIL>
 "00110000000000000000000000000001", -- 293 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 294 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 295 PROG #<NUMBER 2>
 "00000000010010011000000100100111", -- 296 PROG #<CONS 294 295>
 "00110000000000000000000000001101", -- 297 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 298 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 299 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 300 PROG #<NUMBER 1>
 "00000000010010101100000100101100", -- 301 PROG #<CONS 299 300>
 "00110000000000000000000000001101", -- 302 PROG #<NUMBER 13>
 "00110000000000000000000000000010", -- 303 PROG #<NUMBER 2>
 "00110000000000000000000000000001", -- 304 PROG #<NUMBER 1>
 "00110000000000000000000000001101", -- 305 PROG #<NUMBER 13>
 "00110000000000000000000000000010", -- 306 PROG #<NUMBER 2>
 "00110000000000000000000000000001", -- 307 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 308 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 309 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 310 PROG #<NUMBER 0>
 "00000000010011010100000100110110", -- 311 PROG #<CONS 309 310>
 "00110000000000000000000000001111", -- 312 PROG #<NUMBER 15>
 "00110000000000000000000000001101", -- 313 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 314 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 315 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 316 PROG #<NUMBER 1>
 "00000000010011101100000100111100", -- 317 PROG #<CONS 315 316>
 "00110000000000000000000000000100", -- 318 PROG #<NUMBER 4>
 "00110000000000000000000000001001", -- 319 PROG #<NUMBER 9>
 "00000000010011111100000000000000", -- 320 PROG #<CONS 319 0>
 "00000000010011111000000101000000", -- 321 PROG #<CONS 318 320>
 "00000000010011110100000101000001", -- 322 PROG #<CONS 317 321>
 "00000000010011101000000101000010", -- 323 PROG #<CONS 314 322>
 "00000000010011100100000101000011", -- 324 PROG #<CONS 313 323>
 "00000000010011100000000101000100", -- 325 PROG #<CONS 312 324>
 "00000000010011011100000101000101", -- 326 PROG #<CONS 311 325>
 "00000000010011010000000101000110", -- 327 PROG #<CONS 308 326>
 "00000000010011001100000101000111", -- 328 PROG #<CONS 307 327>
 "00000000010011001000000101001000", -- 329 PROG #<CONS 306 328>
 "00000000010011000100000101001001", -- 330 PROG #<CONS 305 329>
 "00000000010011000000000101001010", -- 331 PROG #<CONS 304 330>
 "00000000010010111100000101001011", -- 332 PROG #<CONS 303 331>
 "00000000010010111000000101001100", -- 333 PROG #<CONS 302 332>
 "00000000010010110100000101001101", -- 334 PROG #<CONS 301 333>
 "00000000010010101000000101001110", -- 335 PROG #<CONS 298 334>
 "00000000010010100100000101001111", -- 336 PROG #<CONS 297 335>
 "00000000010010100000000101010000", -- 337 PROG #<CONS 296 336>
 "00000000010010010100000101010001", -- 338 PROG #<CONS 293 337>
 "00000000010010010000000101010010", -- 339 PROG #<CONS 292 338>
 "00000000010010001100000101010011", -- 340 PROG #<CONS 291 339>
 "00110000000000000000000000000101", -- 341 PROG #<NUMBER 5>
 "00000000010101010100000000000000", -- 342 PROG #<CONS 341 0>
 "00000000010101010000000101010110", -- 343 PROG #<CONS 340 342>
 "00000000010010001000000101010111", -- 344 PROG #<CONS 290 343>
 "00000000010001101000000101011000", -- 345 PROG #<CONS 282 344>
 "00000000010001100100000101011001", -- 346 PROG #<CONS 281 345>
 "00000000010001100000000101011010", -- 347 PROG #<CONS 280 346>
 "00000000010001010100000101011011", -- 348 PROG #<CONS 277 347>
 "00000000010001010000000101011100", -- 349 PROG #<CONS 276 348>
 "00000000010001000100000101011101", -- 350 PROG #<CONS 273 349>
 "00110000000000000000000000001101", -- 351 PROG #<NUMBER 13>
 "00110000000000000000000000000011", -- 352 PROG #<NUMBER 3>
 "00110000000000000000000000000010", -- 353 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 354 PROG #<SYMBOL NIL>
 "00110000000000000000000000000001", -- 355 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 356 PROG #<NUMBER 0>
 "00110000000000000000000000000011", -- 357 PROG #<NUMBER 3>
 "00000000010110010000000101100101", -- 358 PROG #<CONS 356 357>
 "00110000000000000000000000001101", -- 359 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 360 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 361 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 362 PROG #<NUMBER 1>
 "00000000010110100100000101101010", -- 363 PROG #<CONS 361 362>
 "00110000000000000000000000001101", -- 364 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 365 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 366 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 367 PROG #<NUMBER 0>
 "00000000010110111000000101101111", -- 368 PROG #<CONS 366 367>
 "00110000000000000000000000001101", -- 369 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 370 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 371 PROG #<NUMBER 1>
 "00110000000000000000000000000101", -- 372 PROG #<NUMBER 5>
 "00000000010111001100000101110100", -- 373 PROG #<CONS 371 372>
 "00110000000000000000000000000100", -- 374 PROG #<NUMBER 4>
 "00110000000000000000000000001000", -- 375 PROG #<NUMBER 8>
 "00110000000000000000000000000010", -- 376 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 377 PROG #<SYMBOL NIL>
 "00110000000000000000000000001001", -- 378 PROG #<NUMBER 9>
 "00000000010111101000000000000000", -- 379 PROG #<CONS 378 0>
 "00000000010111100100000101111011", -- 380 PROG #<CONS 377 379>
 "00000000010111100000000101111100", -- 381 PROG #<CONS 376 380>
 "00110000000000000000000000000010", -- 382 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 383 PROG #<SYMBOL NIL>
 "00110000000000000000000000000001", -- 384 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 385 PROG #<NUMBER 0>
 "00110000000000000000000000000011", -- 386 PROG #<NUMBER 3>
 "00000000011000000100000110000010", -- 387 PROG #<CONS 385 386>
 "00110000000000000000000000000001", -- 388 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 389 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 390 PROG #<NUMBER 1>
 "00000000011000010100000110000110", -- 391 PROG #<CONS 389 390>
 "00110000000000000000000000000001", -- 392 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 393 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 394 PROG #<NUMBER 0>
 "00000000011000100100000110001010", -- 395 PROG #<CONS 393 394>
 "00110000000000000000000000001101", -- 396 PROG #<NUMBER 13>
 "00110000000000000000000000001101", -- 397 PROG #<NUMBER 13>
 "00110000000000000000000000001101", -- 398 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 399 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 400 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 401 PROG #<NUMBER 2>
 "00000000011001000000000110010001", -- 402 PROG #<CONS 400 401>
 "00110000000000000000000000001101", -- 403 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 404 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 405 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 406 PROG #<NUMBER 0>
 "00000000011001010100000110010110", -- 407 PROG #<CONS 405 406>
 "00110000000000000000000000001101", -- 408 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 409 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 410 PROG #<NUMBER 1>
 "00110000000000000000000000000100", -- 411 PROG #<NUMBER 4>
 "00000000011001101000000110011011", -- 412 PROG #<CONS 410 411>
 "00110000000000000000000000000100", -- 413 PROG #<NUMBER 4>
 "00110000000000000000000000001001", -- 414 PROG #<NUMBER 9>
 "00000000011001111000000000000000", -- 415 PROG #<CONS 414 0>
 "00000000011001110100000110011111", -- 416 PROG #<CONS 413 415>
 "00000000011001110000000110100000", -- 417 PROG #<CONS 412 416>
 "00000000011001100100000110100001", -- 418 PROG #<CONS 409 417>
 "00000000011001100000000110100010", -- 419 PROG #<CONS 408 418>
 "00000000011001011100000110100011", -- 420 PROG #<CONS 407 419>
 "00000000011001010000000110100100", -- 421 PROG #<CONS 404 420>
 "00000000011001001100000110100101", -- 422 PROG #<CONS 403 421>
 "00000000011001001000000110100110", -- 423 PROG #<CONS 402 422>
 "00000000011000111100000110100111", -- 424 PROG #<CONS 399 423>
 "00000000011000111000000110101000", -- 425 PROG #<CONS 398 424>
 "00000000011000110100000110101001", -- 426 PROG #<CONS 397 425>
 "00000000011000110000000110101010", -- 427 PROG #<CONS 396 426>
 "00000000011000101100000110101011", -- 428 PROG #<CONS 395 427>
 "00000000011000100000000110101100", -- 429 PROG #<CONS 392 428>
 "00000000011000011100000110101101", -- 430 PROG #<CONS 391 429>
 "00000000011000010000000110101110", -- 431 PROG #<CONS 388 430>
 "00000000011000001100000110101111", -- 432 PROG #<CONS 387 431>
 "00000000011000000000000110110000", -- 433 PROG #<CONS 384 432>
 "00000000010111111100000110110001", -- 434 PROG #<CONS 383 433>
 "00000000010111111000000110110010", -- 435 PROG #<CONS 382 434>
 "00110000000000000000000000000101", -- 436 PROG #<NUMBER 5>
 "00000000011011010000000000000000", -- 437 PROG #<CONS 436 0>
 "00000000011011001100000110110101", -- 438 PROG #<CONS 435 437>
 "00000000010111110100000110110110", -- 439 PROG #<CONS 381 438>
 "00000000010111011100000110110111", -- 440 PROG #<CONS 375 439>
 "00000000010111011000000110111000", -- 441 PROG #<CONS 374 440>
 "00000000010111010100000110111001", -- 442 PROG #<CONS 373 441>
 "00000000010111001000000110111010", -- 443 PROG #<CONS 370 442>
 "00000000010111000100000110111011", -- 444 PROG #<CONS 369 443>
 "00000000010111000000000110111100", -- 445 PROG #<CONS 368 444>
 "00000000010110110100000110111101", -- 446 PROG #<CONS 365 445>
 "00000000010110110000000110111110", -- 447 PROG #<CONS 364 446>
 "00000000010110101100000110111111", -- 448 PROG #<CONS 363 447>
 "00000000010110100000000111000000", -- 449 PROG #<CONS 360 448>
 "00000000010110011100000111000001", -- 450 PROG #<CONS 359 449>
 "00000000010110011000000111000010", -- 451 PROG #<CONS 358 450>
 "00000000010110001100000111000011", -- 452 PROG #<CONS 355 451>
 "00000000010110001000000111000100", -- 453 PROG #<CONS 354 452>
 "00000000010110000100000111000101", -- 454 PROG #<CONS 353 453>
 "00110000000000000000000000001101", -- 455 PROG #<NUMBER 13>
 "00110000000000000000000000000011", -- 456 PROG #<NUMBER 3>
 "00110000000000000000000000000001", -- 457 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 458 PROG #<NUMBER 0>
 "00110000000000000000000000000100", -- 459 PROG #<NUMBER 4>
 "00000000011100101000000111001011", -- 460 PROG #<CONS 458 459>
 "00110000000000000000000000000010", -- 461 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 462 PROG #<SYMBOL NIL>
 "00110000000000000000000000001110", -- 463 PROG #<NUMBER 14>
 "00110000000000000000000000001000", -- 464 PROG #<NUMBER 8>
 "00110000000000000000000000000001", -- 465 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 466 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 467 PROG #<NUMBER 1>
 "00000000011101001000000111010011", -- 468 PROG #<CONS 466 467>
 "00110000000000000000000000000001", -- 469 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 470 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 471 PROG #<NUMBER 2>
 "00000000011101011000000111010111", -- 472 PROG #<CONS 470 471>
 "00110000000000000000000000001110", -- 473 PROG #<NUMBER 14>
 "00110000000000000000000000001000", -- 474 PROG #<NUMBER 8>
 "00110000000000000000000000000010", -- 475 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 476 PROG #<SYMBOL NIL>
 "00110000000000000000000000001001", -- 477 PROG #<NUMBER 9>
 "00000000011101110100000000000000", -- 478 PROG #<CONS 477 0>
 "00000000011101110000000111011110", -- 479 PROG #<CONS 476 478>
 "00000000011101101100000111011111", -- 480 PROG #<CONS 475 479>
 "00110000000000000000000000000010", -- 481 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 482 PROG #<SYMBOL NIL>
 "00110000000000000000000000000001", -- 483 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 484 PROG #<NUMBER 0>
 "00110000000000000000000000000011", -- 485 PROG #<NUMBER 3>
 "00000000011110010000000111100101", -- 486 PROG #<CONS 484 485>
 "00110000000000000000000000001101", -- 487 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 488 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 489 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 490 PROG #<NUMBER 2>
 "00000000011110100100000111101010", -- 491 PROG #<CONS 489 490>
 "00110000000000000000000000001101", -- 492 PROG #<NUMBER 13>
 "00110000000000000000000000000010", -- 493 PROG #<NUMBER 2>
 "00110000000000000000000000000001", -- 494 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 495 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 496 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 497 PROG #<NUMBER 1>
 "00000000011111000000000111110001", -- 498 PROG #<CONS 496 497>
 "00110000000000000000000000001111", -- 499 PROG #<NUMBER 15>
 "00110000000000000000000000001101", -- 500 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 501 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 502 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 503 PROG #<NUMBER 0>
 "00000000011111011000000111110111", -- 504 PROG #<CONS 502 503>
 "00110000000000000000000000001101", -- 505 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 506 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 507 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 508 PROG #<NUMBER 1>
 "00000000011111101100000111111100", -- 509 PROG #<CONS 507 508>
 "00110000000000000000000000000100", -- 510 PROG #<NUMBER 4>
 "00110000000000000000000000001001", -- 511 PROG #<NUMBER 9>
 "00000000011111111100000000000000", -- 512 PROG #<CONS 511 0>
 "00000000011111111000001000000000", -- 513 PROG #<CONS 510 512>
 "00000000011111110100001000000001", -- 514 PROG #<CONS 509 513>
 "00000000011111101000001000000010", -- 515 PROG #<CONS 506 514>
 "00000000011111100100001000000011", -- 516 PROG #<CONS 505 515>
 "00000000011111100000001000000100", -- 517 PROG #<CONS 504 516>
 "00000000011111010100001000000101", -- 518 PROG #<CONS 501 517>
 "00000000011111010000001000000110", -- 519 PROG #<CONS 500 518>
 "00000000011111001100001000000111", -- 520 PROG #<CONS 499 519>
 "00000000011111001000001000001000", -- 521 PROG #<CONS 498 520>
 "00000000011110111100001000001001", -- 522 PROG #<CONS 495 521>
 "00000000011110111000001000001010", -- 523 PROG #<CONS 494 522>
 "00000000011110110100001000001011", -- 524 PROG #<CONS 493 523>
 "00000000011110110000001000001100", -- 525 PROG #<CONS 492 524>
 "00000000011110101100001000001101", -- 526 PROG #<CONS 491 525>
 "00000000011110100000001000001110", -- 527 PROG #<CONS 488 526>
 "00000000011110011100001000001111", -- 528 PROG #<CONS 487 527>
 "00000000011110011000001000010000", -- 529 PROG #<CONS 486 528>
 "00000000011110001100001000010001", -- 530 PROG #<CONS 483 529>
 "00000000011110001000001000010010", -- 531 PROG #<CONS 482 530>
 "00000000011110000100001000010011", -- 532 PROG #<CONS 481 531>
 "00110000000000000000000000001001", -- 533 PROG #<NUMBER 9>
 "00000000100001010100000000000000", -- 534 PROG #<CONS 533 0>
 "00000000100001010000001000010110", -- 535 PROG #<CONS 532 534>
 "00000000011110000000001000010111", -- 536 PROG #<CONS 480 535>
 "00000000011101101000001000011000", -- 537 PROG #<CONS 474 536>
 "00000000011101100100001000011001", -- 538 PROG #<CONS 473 537>
 "00000000011101100000001000011010", -- 539 PROG #<CONS 472 538>
 "00000000011101010100001000011011", -- 540 PROG #<CONS 469 539>
 "00000000011101010000001000011100", -- 541 PROG #<CONS 468 540>
 "00000000011101000100001000011101", -- 542 PROG #<CONS 465 541>
 "00110000000000000000000000000001", -- 543 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 544 PROG #<NUMBER 0>
 "00110000000000000000000000000100", -- 545 PROG #<NUMBER 4>
 "00000000100010000000001000100001", -- 546 PROG #<CONS 544 545>
 "00110000000000000000000000001001", -- 547 PROG #<NUMBER 9>
 "00000000100010001100000000000000", -- 548 PROG #<CONS 547 0>
 "00000000100010001000001000100100", -- 549 PROG #<CONS 546 548>
 "00000000100001111100001000100101", -- 550 PROG #<CONS 543 549>
 "00110000000000000000000000000101", -- 551 PROG #<NUMBER 5>
 "00000000100010011100000000000000", -- 552 PROG #<CONS 551 0>
 "00000000100010011000001000101000", -- 553 PROG #<CONS 550 552>
 "00000000100001111000001000101001", -- 554 PROG #<CONS 542 553>
 "00000000011101000000001000101010", -- 555 PROG #<CONS 464 554>
 "00000000011100111100001000101011", -- 556 PROG #<CONS 463 555>
 "00000000011100111000001000101100", -- 557 PROG #<CONS 462 556>
 "00000000011100110100001000101101", -- 558 PROG #<CONS 461 557>
 "00000000011100110000001000101110", -- 559 PROG #<CONS 460 558>
 "00000000011100100100001000101111", -- 560 PROG #<CONS 457 559>
 "00110000000000000000000000001101", -- 561 PROG #<NUMBER 13>
 "00110000000000000000000000000011", -- 562 PROG #<NUMBER 3>
 "00110000000000000000000000000010", -- 563 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 564 PROG #<SYMBOL NIL>
 "00110000000000000000000000000010", -- 565 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 566 PROG #<SYMBOL NIL>
 "00110000000000000000000000000001", -- 567 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 568 PROG #<NUMBER 0>
 "00110000000000000000000000000011", -- 569 PROG #<NUMBER 3>
 "00000000100011100000001000111001", -- 570 PROG #<CONS 568 569>
 "00110000000000000000000000001101", -- 571 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 572 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 573 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 574 PROG #<NUMBER 2>
 "00000000100011110100001000111110", -- 575 PROG #<CONS 573 574>
 "00110000000000000000000000001101", -- 576 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 577 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 578 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 579 PROG #<NUMBER 1>
 "00000000100100001000001001000011", -- 580 PROG #<CONS 578 579>
 "00110000000000000000000000001101", -- 581 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 582 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 583 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 584 PROG #<NUMBER 0>
 "00000000100100011100001001001000", -- 585 PROG #<CONS 583 584>
 "00110000000000000000000000001101", -- 586 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 587 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 588 PROG #<NUMBER 1>
 "00110000000000000000000000000011", -- 589 PROG #<NUMBER 3>
 "00000000100100110000001001001101", -- 590 PROG #<CONS 588 589>
 "00110000000000000000000000000100", -- 591 PROG #<NUMBER 4>
 "00110000000000000000000000001101", -- 592 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 593 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 594 PROG #<NUMBER 0>
 "00110000000000000000000000000011", -- 595 PROG #<NUMBER 3>
 "00000000100101001000001001010011", -- 596 PROG #<CONS 594 595>
 "00110000000000000000000000001101", -- 597 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 598 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 599 PROG #<NUMBER 0>
 "00110000000000000000000000000010", -- 600 PROG #<NUMBER 2>
 "00000000100101011100001001011000", -- 601 PROG #<CONS 599 600>
 "00110000000000000000000000001101", -- 602 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 603 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 604 PROG #<NUMBER 0>
 "00110000000000000000000000000001", -- 605 PROG #<NUMBER 1>
 "00000000100101110000001001011101", -- 606 PROG #<CONS 604 605>
 "00110000000000000000000000001101", -- 607 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 608 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 609 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 610 PROG #<NUMBER 0>
 "00000000100110000100001001100010", -- 611 PROG #<CONS 609 610>
 "00110000000000000000000000001101", -- 612 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 613 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 614 PROG #<NUMBER 1>
 "00110000000000000000000000000010", -- 615 PROG #<NUMBER 2>
 "00000000100110011000001001100111", -- 616 PROG #<CONS 614 615>
 "00110000000000000000000000000100", -- 617 PROG #<NUMBER 4>
 "00110000000000000000000000000101", -- 618 PROG #<NUMBER 5>
 "00000000100110101000000000000000", -- 619 PROG #<CONS 618 0>
 "00000000100110100100001001101011", -- 620 PROG #<CONS 617 619>
 "00000000100110100000001001101100", -- 621 PROG #<CONS 616 620>
 "00000000100110010100001001101101", -- 622 PROG #<CONS 613 621>
 "00000000100110010000001001101110", -- 623 PROG #<CONS 612 622>
 "00000000100110001100001001101111", -- 624 PROG #<CONS 611 623>
 "00000000100110000000001001110000", -- 625 PROG #<CONS 608 624>
 "00000000100101111100001001110001", -- 626 PROG #<CONS 607 625>
 "00000000100101111000001001110010", -- 627 PROG #<CONS 606 626>
 "00000000100101101100001001110011", -- 628 PROG #<CONS 603 627>
 "00000000100101101000001001110100", -- 629 PROG #<CONS 602 628>
 "00000000100101100100001001110101", -- 630 PROG #<CONS 601 629>
 "00000000100101011000001001110110", -- 631 PROG #<CONS 598 630>
 "00000000100101010100001001110111", -- 632 PROG #<CONS 597 631>
 "00000000100101010000001001111000", -- 633 PROG #<CONS 596 632>
 "00000000100101000100001001111001", -- 634 PROG #<CONS 593 633>
 "00000000100101000000001001111010", -- 635 PROG #<CONS 592 634>
 "00000000100100111100001001111011", -- 636 PROG #<CONS 591 635>
 "00000000100100111000001001111100", -- 637 PROG #<CONS 590 636>
 "00000000100100101100001001111101", -- 638 PROG #<CONS 587 637>
 "00000000100100101000001001111110", -- 639 PROG #<CONS 586 638>
 "00000000100100100100001001111111", -- 640 PROG #<CONS 585 639>
 "00000000100100011000001010000000", -- 641 PROG #<CONS 582 640>
 "00000000100100010100001010000001", -- 642 PROG #<CONS 581 641>
 "00000000100100010000001010000010", -- 643 PROG #<CONS 580 642>
 "00000000100100000100001010000011", -- 644 PROG #<CONS 577 643>
 "00000000100100000000001010000100", -- 645 PROG #<CONS 576 644>
 "00000000100011111100001010000101", -- 646 PROG #<CONS 575 645>
 "00000000100011110000001010000110", -- 647 PROG #<CONS 572 646>
 "00000000100011101100001010000111", -- 648 PROG #<CONS 571 647>
 "00000000100011101000001010001000", -- 649 PROG #<CONS 570 648>
 "00000000100011011100001010001001", -- 650 PROG #<CONS 567 649>
 "00000000100011011000001010001010", -- 651 PROG #<CONS 566 650>
 "00000000100011010100001010001011", -- 652 PROG #<CONS 565 651>
 "00000000100011010000001010001100", -- 653 PROG #<CONS 564 652>
 "00000000100011001100001010001101", -- 654 PROG #<CONS 563 653>
 "00110000000000000000000000001101", -- 655 PROG #<NUMBER 13>
 "00110000000000000000000000000011", -- 656 PROG #<NUMBER 3>
 "00110000000000000000000000000010", -- 657 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 658 PROG #<SYMBOL NIL>
 "00110000000000000000000000000010", -- 659 PROG #<NUMBER 2>
 "00100000000000000000000000000000", -- 660 PROG #<SYMBOL NIL>
 "00110000000000000000000000001101", -- 661 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 662 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 663 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 664 PROG #<NUMBER 0>
 "00000000101001011100001010011000", -- 665 PROG #<CONS 663 664>
 "00110000000000000000000000001101", -- 666 PROG #<NUMBER 13>
 "00110000000000000000000000000010", -- 667 PROG #<NUMBER 2>
 "00110000000000000000000000000001", -- 668 PROG #<NUMBER 1>
 "00110000000000000000000000001101", -- 669 PROG #<NUMBER 13>
 "00110000000000000000000000000010", -- 670 PROG #<NUMBER 2>
 "00110000000000000000000000000001", -- 671 PROG #<NUMBER 1>
 "00110000000000000000000000001101", -- 672 PROG #<NUMBER 13>
 "00110000000000000000000000000001", -- 673 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 674 PROG #<NUMBER 1>
 "00110000000000000000000000000001", -- 675 PROG #<NUMBER 1>
 "00000000101010001000001010100011", -- 676 PROG #<CONS 674 675>
 "00110000000000000000000000000100", -- 677 PROG #<NUMBER 4>
 "00110000000000000000000000000101", -- 678 PROG #<NUMBER 5>
 "00000000101010011000000000000000", -- 679 PROG #<CONS 678 0>
 "00000000101010010100001010100111", -- 680 PROG #<CONS 677 679>
 "00000000101010010000001010101000", -- 681 PROG #<CONS 676 680>
 "00000000101010000100001010101001", -- 682 PROG #<CONS 673 681>
 "00000000101010000000001010101010", -- 683 PROG #<CONS 672 682>
 "00000000101001111100001010101011", -- 684 PROG #<CONS 671 683>
 "00000000101001111000001010101100", -- 685 PROG #<CONS 670 684>
 "00000000101001110100001010101101", -- 686 PROG #<CONS 669 685>
 "00000000101001110000001010101110", -- 687 PROG #<CONS 668 686>
 "00000000101001101100001010101111", -- 688 PROG #<CONS 667 687>
 "00000000101001101000001010110000", -- 689 PROG #<CONS 666 688>
 "00000000101001100100001010110001", -- 690 PROG #<CONS 665 689>
 "00000000101001011000001010110010", -- 691 PROG #<CONS 662 690>
 "00000000101001010100001010110011", -- 692 PROG #<CONS 661 691>
 "00000000101001010000001010110100", -- 693 PROG #<CONS 660 692>
 "00000000101001001100001010110101", -- 694 PROG #<CONS 659 693>
 "00000000101001001000001010110110", -- 695 PROG #<CONS 658 694>
 "00000000101001000100001010110111", -- 696 PROG #<CONS 657 695>
 "00110000000000000000000000001101", -- 697 PROG #<NUMBER 13>
 "00110000000000000000000000000011", -- 698 PROG #<NUMBER 3>
 "00110000000000000000000000000001", -- 699 PROG #<NUMBER 1>
 "00110000000000000000000000000000", -- 700 PROG #<NUMBER 0>
 "00110000000000000000000000000000", -- 701 PROG #<NUMBER 0>
 "00000000101011110000001010111101", -- 702 PROG #<CONS 700 701>
 "00110000000000000000000000000101", -- 703 PROG #<NUMBER 5>
 "00000000101011111100000000000000", -- 704 PROG #<CONS 703 0>
 "00000000101011111000001011000000", -- 705 PROG #<CONS 702 704>
 "00000000101011101100001011000001", -- 706 PROG #<CONS 699 705>
 "00110000000000000000000000000111", -- 707 PROG #<NUMBER 7>
 "00110000000000000000000000000100", -- 708 PROG #<NUMBER 4>
 "00110000000000000000000000010101", -- 709 PROG #<NUMBER 21>
 "00000000101100010100000000000000", -- 710 PROG #<CONS 709 0>
 "00000000101100010000001011000110", -- 711 PROG #<CONS 708 710>
 "00000000101100001100001011000111", -- 712 PROG #<CONS 707 711>
 "00000000101100001000001011001000", -- 713 PROG #<CONS 706 712>
 "00000000101011101000001011001001", -- 714 PROG #<CONS 698 713>
 "00000000101011100100001011001010", -- 715 PROG #<CONS 697 714>
 "00000000101011100000001011001011", -- 716 PROG #<CONS 696 715>
 "00000000101001000000001011001100", -- 717 PROG #<CONS 656 716>
 "00000000101000111100001011001101", -- 718 PROG #<CONS 655 717>
 "00000000101000111000001011001110", -- 719 PROG #<CONS 654 718>
 "00000000100011001000001011001111", -- 720 PROG #<CONS 562 719>
 "00000000100011000100001011010000", -- 721 PROG #<CONS 561 720>
 "00000000100011000000001011010001", -- 722 PROG #<CONS 560 721>
 "00000000011100100000001011010010", -- 723 PROG #<CONS 456 722>
 "00000000011100011100001011010011", -- 724 PROG #<CONS 455 723>
 "00000000011100011000001011010100", -- 725 PROG #<CONS 454 724>
 "00000000010110000000001011010101", -- 726 PROG #<CONS 352 725>
 "00000000010101111100001011010110", -- 727 PROG #<CONS 351 726>
 "00000000010101111000001011010111", -- 728 PROG #<CONS 350 727>
 "00000000010001000000001011011000", -- 729 PROG #<CONS 272 728>
 "00000000010000111100001011011001", -- 730 PROG #<CONS 271 729>
 "00000000010000111000001011011010", -- 731 PROG #<CONS 270 730>
 "00000000001011100000001011011011", -- 732 PROG #<CONS 184 731>
 "00000000001011011100001011011100", -- 733 PROG #<CONS 183 732>
 "00000000001011011000001011011101", -- 734 PROG #<CONS 182 733>
 "00000000000000011000001011011110", -- 735 PROG #<CONS 6 734>
 "00000000000000010100001011011111", -- 736 PROG #<CONS 5 735>
 "00000000000000010000001011100000", -- 737 PROG #<CONS 4 736>
 "00000000000000001100001011100001", -- 738 PROG #<CONS 3 737>
 "00110000000000000000000000001011", -- 739 ARG #<NUMBER 11>
 "00000000101110001100000000000000", -- 740 ARG #<CONS 739 0>
 "00000000101110010000000000000000", -- 741 ARG #<CONS 740 0>
 "00000000101110001000001011100101", -- 742 PROBLEM #<CONS 738 741>
 "00000000000000000000001011101000", -- 743 FREE #<CONS 0 744>
 "00000000000000000000001011101001", -- 744 FREE #<CONS 0 745>
 "00000000000000000000001011101010", -- 745 FREE #<CONS 0 746>
 "00000000000000000000001011101011", -- 746 FREE #<CONS 0 747>
 "00000000000000000000001011101100", -- 747 FREE #<CONS 0 748>
 "00000000000000000000001011101101", -- 748 FREE #<CONS 0 749>
 "00000000000000000000001011101110", -- 749 FREE #<CONS 0 750>
 "00000000000000000000001011101111", -- 750 FREE #<CONS 0 751>
 "00000000000000000000001011110000", -- 751 FREE #<CONS 0 752>
 "00000000000000000000001011110001", -- 752 FREE #<CONS 0 753>
 "00000000000000000000001011110010", -- 753 FREE #<CONS 0 754>
 "00000000000000000000001011110011", -- 754 FREE #<CONS 0 755>
 "00000000000000000000001011110100", -- 755 FREE #<CONS 0 756>
 "00000000000000000000001011110101", -- 756 FREE #<CONS 0 757>
 "00000000000000000000001011110110", -- 757 FREE #<CONS 0 758>
 "00000000000000000000001011110111", -- 758 FREE #<CONS 0 759>
 "00000000000000000000001011111000", -- 759 FREE #<CONS 0 760>
 "00000000000000000000001011111001", -- 760 FREE #<CONS 0 761>
 "00000000000000000000001011111010", -- 761 FREE #<CONS 0 762>
 "00000000000000000000001011111011", -- 762 FREE #<CONS 0 763>
 "00000000000000000000001011111100", -- 763 FREE #<CONS 0 764>
 "00000000000000000000001011111101", -- 764 FREE #<CONS 0 765>
 "00000000000000000000001011111110", -- 765 FREE #<CONS 0 766>
 "00000000000000000000001011111111", -- 766 FREE #<CONS 0 767>
 "00000000000000000000001100000000", -- 767 FREE #<CONS 0 768>
 "00000000000000000000001100000001", -- 768 FREE #<CONS 0 769>
 "00000000000000000000001100000010", -- 769 FREE #<CONS 0 770>
 "00000000000000000000001100000011", -- 770 FREE #<CONS 0 771>
 "00000000000000000000001100000100", -- 771 FREE #<CONS 0 772>
 "00000000000000000000001100000101", -- 772 FREE #<CONS 0 773>
 "00000000000000000000001100000110", -- 773 FREE #<CONS 0 774>
 "00000000000000000000001100000111", -- 774 FREE #<CONS 0 775>
 "00000000000000000000001100001000", -- 775 FREE #<CONS 0 776>
 "00000000000000000000001100001001", -- 776 FREE #<CONS 0 777>
 "00000000000000000000001100001010", -- 777 FREE #<CONS 0 778>
 "00000000000000000000001100001011", -- 778 FREE #<CONS 0 779>
 "00000000000000000000001100001100", -- 779 FREE #<CONS 0 780>
 "00000000000000000000001100001101", -- 780 FREE #<CONS 0 781>
 "00000000000000000000001100001110", -- 781 FREE #<CONS 0 782>
 "00000000000000000000001100001111", -- 782 FREE #<CONS 0 783>
 "00000000000000000000001100010000", -- 783 FREE #<CONS 0 784>
 "00000000000000000000001100010001", -- 784 FREE #<CONS 0 785>
 "00000000000000000000001100010010", -- 785 FREE #<CONS 0 786>
 "00000000000000000000001100010011", -- 786 FREE #<CONS 0 787>
 "00000000000000000000001100010100", -- 787 FREE #<CONS 0 788>
 "00000000000000000000001100010101", -- 788 FREE #<CONS 0 789>
 "00000000000000000000001100010110", -- 789 FREE #<CONS 0 790>
 "00000000000000000000001100010111", -- 790 FREE #<CONS 0 791>
 "00000000000000000000001100011000", -- 791 FREE #<CONS 0 792>
 "00000000000000000000001100011001", -- 792 FREE #<CONS 0 793>
 "00000000000000000000001100011010", -- 793 FREE #<CONS 0 794>
 "00000000000000000000001100011011", -- 794 FREE #<CONS 0 795>
 "00000000000000000000001100011100", -- 795 FREE #<CONS 0 796>
 "00000000000000000000001100011101", -- 796 FREE #<CONS 0 797>
 "00000000000000000000001100011110", -- 797 FREE #<CONS 0 798>
 "00000000000000000000001100011111", -- 798 FREE #<CONS 0 799>
 "00000000000000000000001100100000", -- 799 FREE #<CONS 0 800>
 "00000000000000000000001100100001", -- 800 FREE #<CONS 0 801>
 "00000000000000000000001100100010", -- 801 FREE #<CONS 0 802>
 "00000000000000000000001100100011", -- 802 FREE #<CONS 0 803>
 "00000000000000000000001100100100", -- 803 FREE #<CONS 0 804>
 "00000000000000000000001100100101", -- 804 FREE #<CONS 0 805>
 "00000000000000000000001100100110", -- 805 FREE #<CONS 0 806>
 "00000000000000000000001100100111", -- 806 FREE #<CONS 0 807>
 "00000000000000000000001100101000", -- 807 FREE #<CONS 0 808>
 "00000000000000000000001100101001", -- 808 FREE #<CONS 0 809>
 "00000000000000000000001100101010", -- 809 FREE #<CONS 0 810>
 "00000000000000000000001100101011", -- 810 FREE #<CONS 0 811>
 "00000000000000000000001100101100", -- 811 FREE #<CONS 0 812>
 "00000000000000000000001100101101", -- 812 FREE #<CONS 0 813>
 "00000000000000000000001100101110", -- 813 FREE #<CONS 0 814>
 "00000000000000000000001100101111", -- 814 FREE #<CONS 0 815>
 "00000000000000000000001100110000", -- 815 FREE #<CONS 0 816>
 "00000000000000000000001100110001", -- 816 FREE #<CONS 0 817>
 "00000000000000000000001100110010", -- 817 FREE #<CONS 0 818>
 "00000000000000000000001100110011", -- 818 FREE #<CONS 0 819>
 "00000000000000000000001100110100", -- 819 FREE #<CONS 0 820>
 "00000000000000000000001100110101", -- 820 FREE #<CONS 0 821>
 "00000000000000000000001100110110", -- 821 FREE #<CONS 0 822>
 "00000000000000000000001100110111", -- 822 FREE #<CONS 0 823>
 "00000000000000000000001100111000", -- 823 FREE #<CONS 0 824>
 "00000000000000000000001100111001", -- 824 FREE #<CONS 0 825>
 "00000000000000000000001100111010", -- 825 FREE #<CONS 0 826>
 "00000000000000000000001100111011", -- 826 FREE #<CONS 0 827>
 "00000000000000000000001100111100", -- 827 FREE #<CONS 0 828>
 "00000000000000000000001100111101", -- 828 FREE #<CONS 0 829>
 "00000000000000000000001100111110", -- 829 FREE #<CONS 0 830>
 "00000000000000000000001100111111", -- 830 FREE #<CONS 0 831>
 "00000000000000000000001101000000", -- 831 FREE #<CONS 0 832>
 "00000000000000000000001101000001", -- 832 FREE #<CONS 0 833>
 "00000000000000000000001101000010", -- 833 FREE #<CONS 0 834>
 "00000000000000000000001101000011", -- 834 FREE #<CONS 0 835>
 "00000000000000000000001101000100", -- 835 FREE #<CONS 0 836>
 "00000000000000000000001101000101", -- 836 FREE #<CONS 0 837>
 "00000000000000000000001101000110", -- 837 FREE #<CONS 0 838>
 "00000000000000000000001101000111", -- 838 FREE #<CONS 0 839>
 "00000000000000000000001101001000", -- 839 FREE #<CONS 0 840>
 "00000000000000000000001101001001", -- 840 FREE #<CONS 0 841>
 "00000000000000000000001101001010", -- 841 FREE #<CONS 0 842>
 "00000000000000000000001101001011", -- 842 FREE #<CONS 0 843>
 "00000000000000000000001101001100", -- 843 FREE #<CONS 0 844>
 "00000000000000000000001101001101", -- 844 FREE #<CONS 0 845>
 "00000000000000000000001101001110", -- 845 FREE #<CONS 0 846>
 "00000000000000000000001101001111", -- 846 FREE #<CONS 0 847>
 "00000000000000000000001101010000", -- 847 FREE #<CONS 0 848>
 "00000000000000000000001101010001", -- 848 FREE #<CONS 0 849>
 "00000000000000000000001101010010", -- 849 FREE #<CONS 0 850>
 "00000000000000000000001101010011", -- 850 FREE #<CONS 0 851>
 "00000000000000000000001101010100", -- 851 FREE #<CONS 0 852>
 "00000000000000000000001101010101", -- 852 FREE #<CONS 0 853>
 "00000000000000000000001101010110", -- 853 FREE #<CONS 0 854>
 "00000000000000000000001101010111", -- 854 FREE #<CONS 0 855>
 "00000000000000000000001101011000", -- 855 FREE #<CONS 0 856>
 "00000000000000000000001101011001", -- 856 FREE #<CONS 0 857>
 "00000000000000000000001101011010", -- 857 FREE #<CONS 0 858>
 "00000000000000000000001101011011", -- 858 FREE #<CONS 0 859>
 "00000000000000000000001101011100", -- 859 FREE #<CONS 0 860>
 "00000000000000000000001101011101", -- 860 FREE #<CONS 0 861>
 "00000000000000000000001101011110", -- 861 FREE #<CONS 0 862>
 "00000000000000000000001101011111", -- 862 FREE #<CONS 0 863>
 "00000000000000000000001101100000", -- 863 FREE #<CONS 0 864>
 "00000000000000000000001101100001", -- 864 FREE #<CONS 0 865>
 "00000000000000000000001101100010", -- 865 FREE #<CONS 0 866>
 "00000000000000000000001101100011", -- 866 FREE #<CONS 0 867>
 "00000000000000000000001101100100", -- 867 FREE #<CONS 0 868>
 "00000000000000000000001101100101", -- 868 FREE #<CONS 0 869>
 "00000000000000000000001101100110", -- 869 FREE #<CONS 0 870>
 "00000000000000000000001101100111", -- 870 FREE #<CONS 0 871>
 "00000000000000000000001101101000", -- 871 FREE #<CONS 0 872>
 "00000000000000000000001101101001", -- 872 FREE #<CONS 0 873>
 "00000000000000000000001101101010", -- 873 FREE #<CONS 0 874>
 "00000000000000000000001101101011", -- 874 FREE #<CONS 0 875>
 "00000000000000000000001101101100", -- 875 FREE #<CONS 0 876>
 "00000000000000000000001101101101", -- 876 FREE #<CONS 0 877>
 "00000000000000000000001101101110", -- 877 FREE #<CONS 0 878>
 "00000000000000000000001101101111", -- 878 FREE #<CONS 0 879>
 "00000000000000000000001101110000", -- 879 FREE #<CONS 0 880>
 "00000000000000000000001101110001", -- 880 FREE #<CONS 0 881>
 "00000000000000000000001101110010", -- 881 FREE #<CONS 0 882>
 "00000000000000000000001101110011", -- 882 FREE #<CONS 0 883>
 "00000000000000000000001101110100", -- 883 FREE #<CONS 0 884>
 "00000000000000000000001101110101", -- 884 FREE #<CONS 0 885>
 "00000000000000000000001101110110", -- 885 FREE #<CONS 0 886>
 "00000000000000000000001101110111", -- 886 FREE #<CONS 0 887>
 "00000000000000000000001101111000", -- 887 FREE #<CONS 0 888>
 "00000000000000000000001101111001", -- 888 FREE #<CONS 0 889>
 "00000000000000000000001101111010", -- 889 FREE #<CONS 0 890>
 "00000000000000000000001101111011", -- 890 FREE #<CONS 0 891>
 "00000000000000000000001101111100", -- 891 FREE #<CONS 0 892>
 "00000000000000000000001101111101", -- 892 FREE #<CONS 0 893>
 "00000000000000000000001101111110", -- 893 FREE #<CONS 0 894>
 "00000000000000000000001101111111", -- 894 FREE #<CONS 0 895>
 "00000000000000000000001110000000", -- 895 FREE #<CONS 0 896>
 "00000000000000000000001110000001", -- 896 FREE #<CONS 0 897>
 "00000000000000000000001110000010", -- 897 FREE #<CONS 0 898>
 "00000000000000000000001110000011", -- 898 FREE #<CONS 0 899>
 "00000000000000000000001110000100", -- 899 FREE #<CONS 0 900>
 "00000000000000000000001110000101", -- 900 FREE #<CONS 0 901>
 "00000000000000000000001110000110", -- 901 FREE #<CONS 0 902>
 "00000000000000000000001110000111", -- 902 FREE #<CONS 0 903>
 "00000000000000000000001110001000", -- 903 FREE #<CONS 0 904>
 "00000000000000000000001110001001", -- 904 FREE #<CONS 0 905>
 "00000000000000000000001110001010", -- 905 FREE #<CONS 0 906>
 "00000000000000000000001110001011", -- 906 FREE #<CONS 0 907>
 "00000000000000000000001110001100", -- 907 FREE #<CONS 0 908>
 "00000000000000000000001110001101", -- 908 FREE #<CONS 0 909>
 "00000000000000000000001110001110", -- 909 FREE #<CONS 0 910>
 "00000000000000000000001110001111", -- 910 FREE #<CONS 0 911>
 "00000000000000000000001110010000", -- 911 FREE #<CONS 0 912>
 "00000000000000000000001110010001", -- 912 FREE #<CONS 0 913>
 "00000000000000000000001110010010", -- 913 FREE #<CONS 0 914>
 "00000000000000000000001110010011", -- 914 FREE #<CONS 0 915>
 "00000000000000000000001110010100", -- 915 FREE #<CONS 0 916>
 "00000000000000000000001110010101", -- 916 FREE #<CONS 0 917>
 "00000000000000000000001110010110", -- 917 FREE #<CONS 0 918>
 "00000000000000000000001110010111", -- 918 FREE #<CONS 0 919>
 "00000000000000000000001110011000", -- 919 FREE #<CONS 0 920>
 "00000000000000000000001110011001", -- 920 FREE #<CONS 0 921>
 "00000000000000000000001110011010", -- 921 FREE #<CONS 0 922>
 "00000000000000000000001110011011", -- 922 FREE #<CONS 0 923>
 "00000000000000000000001110011100", -- 923 FREE #<CONS 0 924>
 "00000000000000000000001110011101", -- 924 FREE #<CONS 0 925>
 "00000000000000000000001110011110", -- 925 FREE #<CONS 0 926>
 "00000000000000000000001110011111", -- 926 FREE #<CONS 0 927>
 "00000000000000000000001110100000", -- 927 FREE #<CONS 0 928>
 "00000000000000000000001110100001", -- 928 FREE #<CONS 0 929>
 "00000000000000000000001110100010", -- 929 FREE #<CONS 0 930>
 "00000000000000000000001110100011", -- 930 FREE #<CONS 0 931>
 "00000000000000000000001110100100", -- 931 FREE #<CONS 0 932>
 "00000000000000000000001110100101", -- 932 FREE #<CONS 0 933>
 "00000000000000000000001110100110", -- 933 FREE #<CONS 0 934>
 "00000000000000000000001110100111", -- 934 FREE #<CONS 0 935>
 "00000000000000000000001110101000", -- 935 FREE #<CONS 0 936>
 "00000000000000000000001110101001", -- 936 FREE #<CONS 0 937>
 "00000000000000000000001110101010", -- 937 FREE #<CONS 0 938>
 "00000000000000000000001110101011", -- 938 FREE #<CONS 0 939>
 "00000000000000000000001110101100", -- 939 FREE #<CONS 0 940>
 "00000000000000000000001110101101", -- 940 FREE #<CONS 0 941>
 "00000000000000000000001110101110", -- 941 FREE #<CONS 0 942>
 "00000000000000000000001110101111", -- 942 FREE #<CONS 0 943>
 "00000000000000000000001110110000", -- 943 FREE #<CONS 0 944>
 "00000000000000000000001110110001", -- 944 FREE #<CONS 0 945>
 "00000000000000000000001110110010", -- 945 FREE #<CONS 0 946>
 "00000000000000000000001110110011", -- 946 FREE #<CONS 0 947>
 "00000000000000000000001110110100", -- 947 FREE #<CONS 0 948>
 "00000000000000000000001110110101", -- 948 FREE #<CONS 0 949>
 "00000000000000000000001110110110", -- 949 FREE #<CONS 0 950>
 "00000000000000000000001110110111", -- 950 FREE #<CONS 0 951>
 "00000000000000000000001110111000", -- 951 FREE #<CONS 0 952>
 "00000000000000000000001110111001", -- 952 FREE #<CONS 0 953>
 "00000000000000000000001110111010", -- 953 FREE #<CONS 0 954>
 "00000000000000000000001110111011", -- 954 FREE #<CONS 0 955>
 "00000000000000000000001110111100", -- 955 FREE #<CONS 0 956>
 "00000000000000000000001110111101", -- 956 FREE #<CONS 0 957>
 "00000000000000000000001110111110", -- 957 FREE #<CONS 0 958>
 "00000000000000000000001110111111", -- 958 FREE #<CONS 0 959>
 "00000000000000000000001111000000", -- 959 FREE #<CONS 0 960>
 "00000000000000000000001111000001", -- 960 FREE #<CONS 0 961>
 "00000000000000000000001111000010", -- 961 FREE #<CONS 0 962>
 "00000000000000000000001111000011", -- 962 FREE #<CONS 0 963>
 "00000000000000000000001111000100", -- 963 FREE #<CONS 0 964>
 "00000000000000000000001111000101", -- 964 FREE #<CONS 0 965>
 "00000000000000000000001111000110", -- 965 FREE #<CONS 0 966>
 "00000000000000000000001111000111", -- 966 FREE #<CONS 0 967>
 "00000000000000000000001111001000", -- 967 FREE #<CONS 0 968>
 "00000000000000000000001111001001", -- 968 FREE #<CONS 0 969>
 "00000000000000000000001111001010", -- 969 FREE #<CONS 0 970>
 "00000000000000000000001111001011", -- 970 FREE #<CONS 0 971>
 "00000000000000000000001111001100", -- 971 FREE #<CONS 0 972>
 "00000000000000000000001111001101", -- 972 FREE #<CONS 0 973>
 "00000000000000000000001111001110", -- 973 FREE #<CONS 0 974>
 "00000000000000000000001111001111", -- 974 FREE #<CONS 0 975>
 "00000000000000000000001111010000", -- 975 FREE #<CONS 0 976>
 "00000000000000000000001111010001", -- 976 FREE #<CONS 0 977>
 "00000000000000000000001111010010", -- 977 FREE #<CONS 0 978>
 "00000000000000000000001111010011", -- 978 FREE #<CONS 0 979>
 "00000000000000000000001111010100", -- 979 FREE #<CONS 0 980>
 "00000000000000000000001111010101", -- 980 FREE #<CONS 0 981>
 "00000000000000000000001111010110", -- 981 FREE #<CONS 0 982>
 "00000000000000000000001111010111", -- 982 FREE #<CONS 0 983>
 "00000000000000000000001111011000", -- 983 FREE #<CONS 0 984>
 "00000000000000000000001111011001", -- 984 FREE #<CONS 0 985>
 "00000000000000000000001111011010", -- 985 FREE #<CONS 0 986>
 "00000000000000000000001111011011", -- 986 FREE #<CONS 0 987>
 "00000000000000000000001111011100", -- 987 FREE #<CONS 0 988>
 "00000000000000000000001111011101", -- 988 FREE #<CONS 0 989>
 "00000000000000000000001111011110", -- 989 FREE #<CONS 0 990>
 "00000000000000000000001111011111", -- 990 FREE #<CONS 0 991>
 "00000000000000000000001111100000", -- 991 FREE #<CONS 0 992>
 "00000000000000000000001111100001", -- 992 FREE #<CONS 0 993>
 "00000000000000000000001111100010", -- 993 FREE #<CONS 0 994>
 "00000000000000000000001111100011", -- 994 FREE #<CONS 0 995>
 "00000000000000000000001111100100", -- 995 FREE #<CONS 0 996>
 "00000000000000000000001111100101", -- 996 FREE #<CONS 0 997>
 "00000000000000000000001111100110", -- 997 FREE #<CONS 0 998>
 "00000000000000000000001111100111", -- 998 FREE #<CONS 0 999>
 "00000000000000000000001111101000", -- 999 FREE #<CONS 0 1000>
 "00000000000000000000001111101001", -- 1000 FREE #<CONS 0 1001>
 "00000000000000000000001111101010", -- 1001 FREE #<CONS 0 1002>
 "00000000000000000000001111101011", -- 1002 FREE #<CONS 0 1003>
 "00000000000000000000001111101100", -- 1003 FREE #<CONS 0 1004>
 "00000000000000000000001111101101", -- 1004 FREE #<CONS 0 1005>
 "00000000000000000000001111101110", -- 1005 FREE #<CONS 0 1006>
 "00000000000000000000001111101111", -- 1006 FREE #<CONS 0 1007>
 "00000000000000000000001111110000", -- 1007 FREE #<CONS 0 1008>
 "00000000000000000000001111110001", -- 1008 FREE #<CONS 0 1009>
 "00000000000000000000001111110010", -- 1009 FREE #<CONS 0 1010>
 "00000000000000000000001111110011", -- 1010 FREE #<CONS 0 1011>
 "00000000000000000000001111110100", -- 1011 FREE #<CONS 0 1012>
 "00000000000000000000001111110101", -- 1012 FREE #<CONS 0 1013>
 "00000000000000000000001111110110", -- 1013 FREE #<CONS 0 1014>
 "00000000000000000000001111110111", -- 1014 FREE #<CONS 0 1015>
 "00000000000000000000001111111000", -- 1015 FREE #<CONS 0 1016>
 "00000000000000000000001111111001", -- 1016 FREE #<CONS 0 1017>
 "00000000000000000000001111111010", -- 1017 FREE #<CONS 0 1018>
 "00000000000000000000001111111011", -- 1018 FREE #<CONS 0 1019>
 "00000000000000000000001111111100", -- 1019 FREE #<CONS 0 1020>
 "00000000000000000000001111111101", -- 1020 FREE #<CONS 0 1021>
 "00000000000000000000001111111110", -- 1021 FREE #<CONS 0 1022>
 "00000000000000000000001111111111", -- 1022 FREE #<CONS 0 1023>
 "00000000000000000000010000000000", -- 1023 FREE #<CONS 0 1024>
 "00000000000000000000010000000001", -- 1024 FREE #<CONS 0 1025>
 "00000000000000000000010000000010", -- 1025 FREE #<CONS 0 1026>
 "00000000000000000000010000000011", -- 1026 FREE #<CONS 0 1027>
 "00000000000000000000010000000100", -- 1027 FREE #<CONS 0 1028>
 "00000000000000000000010000000101", -- 1028 FREE #<CONS 0 1029>
 "00000000000000000000010000000110", -- 1029 FREE #<CONS 0 1030>
 "00000000000000000000010000000111", -- 1030 FREE #<CONS 0 1031>
 "00000000000000000000010000001000", -- 1031 FREE #<CONS 0 1032>
 "00000000000000000000010000001001", -- 1032 FREE #<CONS 0 1033>
 "00000000000000000000010000001010", -- 1033 FREE #<CONS 0 1034>
 "00000000000000000000010000001011", -- 1034 FREE #<CONS 0 1035>
 "00000000000000000000010000001100", -- 1035 FREE #<CONS 0 1036>
 "00000000000000000000010000001101", -- 1036 FREE #<CONS 0 1037>
 "00000000000000000000010000001110", -- 1037 FREE #<CONS 0 1038>
 "00000000000000000000010000001111", -- 1038 FREE #<CONS 0 1039>
 "00000000000000000000010000010000", -- 1039 FREE #<CONS 0 1040>
 "00000000000000000000010000010001", -- 1040 FREE #<CONS 0 1041>
 "00000000000000000000010000010010", -- 1041 FREE #<CONS 0 1042>
 "00000000000000000000010000010011", -- 1042 FREE #<CONS 0 1043>
 "00000000000000000000010000010100", -- 1043 FREE #<CONS 0 1044>
 "00000000000000000000010000010101", -- 1044 FREE #<CONS 0 1045>
 "00000000000000000000010000010110", -- 1045 FREE #<CONS 0 1046>
 "00000000000000000000010000010111", -- 1046 FREE #<CONS 0 1047>
 "00000000000000000000010000011000", -- 1047 FREE #<CONS 0 1048>
 "00000000000000000000010000011001", -- 1048 FREE #<CONS 0 1049>
 "00000000000000000000010000011010", -- 1049 FREE #<CONS 0 1050>
 "00000000000000000000010000011011", -- 1050 FREE #<CONS 0 1051>
 "00000000000000000000010000011100", -- 1051 FREE #<CONS 0 1052>
 "00000000000000000000010000011101", -- 1052 FREE #<CONS 0 1053>
 "00000000000000000000010000011110", -- 1053 FREE #<CONS 0 1054>
 "00000000000000000000010000011111", -- 1054 FREE #<CONS 0 1055>
 "00000000000000000000010000100000", -- 1055 FREE #<CONS 0 1056>
 "00000000000000000000010000100001", -- 1056 FREE #<CONS 0 1057>
 "00000000000000000000010000100010", -- 1057 FREE #<CONS 0 1058>
 "00000000000000000000010000100011", -- 1058 FREE #<CONS 0 1059>
 "00000000000000000000010000100100", -- 1059 FREE #<CONS 0 1060>
 "00000000000000000000010000100101", -- 1060 FREE #<CONS 0 1061>
 "00000000000000000000010000100110", -- 1061 FREE #<CONS 0 1062>
 "00000000000000000000010000100111", -- 1062 FREE #<CONS 0 1063>
 "00000000000000000000010000101000", -- 1063 FREE #<CONS 0 1064>
 "00000000000000000000010000101001", -- 1064 FREE #<CONS 0 1065>
 "00000000000000000000010000101010", -- 1065 FREE #<CONS 0 1066>
 "00000000000000000000010000101011", -- 1066 FREE #<CONS 0 1067>
 "00000000000000000000010000101100", -- 1067 FREE #<CONS 0 1068>
 "00000000000000000000010000101101", -- 1068 FREE #<CONS 0 1069>
 "00000000000000000000010000101110", -- 1069 FREE #<CONS 0 1070>
 "00000000000000000000010000101111", -- 1070 FREE #<CONS 0 1071>
 "00000000000000000000010000110000", -- 1071 FREE #<CONS 0 1072>
 "00000000000000000000010000110001", -- 1072 FREE #<CONS 0 1073>
 "00000000000000000000010000110010", -- 1073 FREE #<CONS 0 1074>
 "00000000000000000000010000110011", -- 1074 FREE #<CONS 0 1075>
 "00000000000000000000010000110100", -- 1075 FREE #<CONS 0 1076>
 "00000000000000000000010000110101", -- 1076 FREE #<CONS 0 1077>
 "00000000000000000000010000110110", -- 1077 FREE #<CONS 0 1078>
 "00000000000000000000010000110111", -- 1078 FREE #<CONS 0 1079>
 "00000000000000000000010000111000", -- 1079 FREE #<CONS 0 1080>
 "00000000000000000000010000111001", -- 1080 FREE #<CONS 0 1081>
 "00000000000000000000010000111010", -- 1081 FREE #<CONS 0 1082>
 "00000000000000000000010000111011", -- 1082 FREE #<CONS 0 1083>
 "00000000000000000000010000111100", -- 1083 FREE #<CONS 0 1084>
 "00000000000000000000010000111101", -- 1084 FREE #<CONS 0 1085>
 "00000000000000000000010000111110", -- 1085 FREE #<CONS 0 1086>
 "00000000000000000000010000111111", -- 1086 FREE #<CONS 0 1087>
 "00000000000000000000010001000000", -- 1087 FREE #<CONS 0 1088>
 "00000000000000000000010001000001", -- 1088 FREE #<CONS 0 1089>
 "00000000000000000000010001000010", -- 1089 FREE #<CONS 0 1090>
 "00000000000000000000010001000011", -- 1090 FREE #<CONS 0 1091>
 "00000000000000000000010001000100", -- 1091 FREE #<CONS 0 1092>
 "00000000000000000000010001000101", -- 1092 FREE #<CONS 0 1093>
 "00000000000000000000010001000110", -- 1093 FREE #<CONS 0 1094>
 "00000000000000000000010001000111", -- 1094 FREE #<CONS 0 1095>
 "00000000000000000000010001001000", -- 1095 FREE #<CONS 0 1096>
 "00000000000000000000010001001001", -- 1096 FREE #<CONS 0 1097>
 "00000000000000000000010001001010", -- 1097 FREE #<CONS 0 1098>
 "00000000000000000000010001001011", -- 1098 FREE #<CONS 0 1099>
 "00000000000000000000010001001100", -- 1099 FREE #<CONS 0 1100>
 "00000000000000000000010001001101", -- 1100 FREE #<CONS 0 1101>
 "00000000000000000000010001001110", -- 1101 FREE #<CONS 0 1102>
 "00000000000000000000010001001111", -- 1102 FREE #<CONS 0 1103>
 "00000000000000000000010001010000", -- 1103 FREE #<CONS 0 1104>
 "00000000000000000000010001010001", -- 1104 FREE #<CONS 0 1105>
 "00000000000000000000010001010010", -- 1105 FREE #<CONS 0 1106>
 "00000000000000000000010001010011", -- 1106 FREE #<CONS 0 1107>
 "00000000000000000000010001010100", -- 1107 FREE #<CONS 0 1108>
 "00000000000000000000010001010101", -- 1108 FREE #<CONS 0 1109>
 "00000000000000000000010001010110", -- 1109 FREE #<CONS 0 1110>
 "00000000000000000000010001010111", -- 1110 FREE #<CONS 0 1111>
 "00000000000000000000010001011000", -- 1111 FREE #<CONS 0 1112>
 "00000000000000000000010001011001", -- 1112 FREE #<CONS 0 1113>
 "00000000000000000000010001011010", -- 1113 FREE #<CONS 0 1114>
 "00000000000000000000010001011011", -- 1114 FREE #<CONS 0 1115>
 "00000000000000000000010001011100", -- 1115 FREE #<CONS 0 1116>
 "00000000000000000000010001011101", -- 1116 FREE #<CONS 0 1117>
 "00000000000000000000010001011110", -- 1117 FREE #<CONS 0 1118>
 "00000000000000000000010001011111", -- 1118 FREE #<CONS 0 1119>
 "00000000000000000000010001100000", -- 1119 FREE #<CONS 0 1120>
 "00000000000000000000010001100001", -- 1120 FREE #<CONS 0 1121>
 "00000000000000000000010001100010", -- 1121 FREE #<CONS 0 1122>
 "00000000000000000000010001100011", -- 1122 FREE #<CONS 0 1123>
 "00000000000000000000010001100100", -- 1123 FREE #<CONS 0 1124>
 "00000000000000000000010001100101", -- 1124 FREE #<CONS 0 1125>
 "00000000000000000000010001100110", -- 1125 FREE #<CONS 0 1126>
 "00000000000000000000010001100111", -- 1126 FREE #<CONS 0 1127>
 "00000000000000000000010001101000", -- 1127 FREE #<CONS 0 1128>
 "00000000000000000000010001101001", -- 1128 FREE #<CONS 0 1129>
 "00000000000000000000010001101010", -- 1129 FREE #<CONS 0 1130>
 "00000000000000000000010001101011", -- 1130 FREE #<CONS 0 1131>
 "00000000000000000000010001101100", -- 1131 FREE #<CONS 0 1132>
 "00000000000000000000010001101101", -- 1132 FREE #<CONS 0 1133>
 "00000000000000000000010001101110", -- 1133 FREE #<CONS 0 1134>
 "00000000000000000000010001101111", -- 1134 FREE #<CONS 0 1135>
 "00000000000000000000010001110000", -- 1135 FREE #<CONS 0 1136>
 "00000000000000000000010001110001", -- 1136 FREE #<CONS 0 1137>
 "00000000000000000000010001110010", -- 1137 FREE #<CONS 0 1138>
 "00000000000000000000010001110011", -- 1138 FREE #<CONS 0 1139>
 "00000000000000000000010001110100", -- 1139 FREE #<CONS 0 1140>
 "00000000000000000000010001110101", -- 1140 FREE #<CONS 0 1141>
 "00000000000000000000010001110110", -- 1141 FREE #<CONS 0 1142>
 "00000000000000000000010001110111", -- 1142 FREE #<CONS 0 1143>
 "00000000000000000000010001111000", -- 1143 FREE #<CONS 0 1144>
 "00000000000000000000010001111001", -- 1144 FREE #<CONS 0 1145>
 "00000000000000000000010001111010", -- 1145 FREE #<CONS 0 1146>
 "00000000000000000000010001111011", -- 1146 FREE #<CONS 0 1147>
 "00000000000000000000010001111100", -- 1147 FREE #<CONS 0 1148>
 "00000000000000000000010001111101", -- 1148 FREE #<CONS 0 1149>
 "00000000000000000000010001111110", -- 1149 FREE #<CONS 0 1150>
 "00000000000000000000010001111111", -- 1150 FREE #<CONS 0 1151>
 "00000000000000000000010010000000", -- 1151 FREE #<CONS 0 1152>
 "00000000000000000000010010000001", -- 1152 FREE #<CONS 0 1153>
 "00000000000000000000010010000010", -- 1153 FREE #<CONS 0 1154>
 "00000000000000000000010010000011", -- 1154 FREE #<CONS 0 1155>
 "00000000000000000000010010000100", -- 1155 FREE #<CONS 0 1156>
 "00000000000000000000010010000101", -- 1156 FREE #<CONS 0 1157>
 "00000000000000000000010010000110", -- 1157 FREE #<CONS 0 1158>
 "00000000000000000000010010000111", -- 1158 FREE #<CONS 0 1159>
 "00000000000000000000010010001000", -- 1159 FREE #<CONS 0 1160>
 "00000000000000000000010010001001", -- 1160 FREE #<CONS 0 1161>
 "00000000000000000000010010001010", -- 1161 FREE #<CONS 0 1162>
 "00000000000000000000010010001011", -- 1162 FREE #<CONS 0 1163>
 "00000000000000000000010010001100", -- 1163 FREE #<CONS 0 1164>
 "00000000000000000000010010001101", -- 1164 FREE #<CONS 0 1165>
 "00000000000000000000010010001110", -- 1165 FREE #<CONS 0 1166>
 "00000000000000000000010010001111", -- 1166 FREE #<CONS 0 1167>
 "00000000000000000000010010010000", -- 1167 FREE #<CONS 0 1168>
 "00000000000000000000010010010001", -- 1168 FREE #<CONS 0 1169>
 "00000000000000000000010010010010", -- 1169 FREE #<CONS 0 1170>
 "00000000000000000000010010010011", -- 1170 FREE #<CONS 0 1171>
 "00000000000000000000010010010100", -- 1171 FREE #<CONS 0 1172>
 "00000000000000000000010010010101", -- 1172 FREE #<CONS 0 1173>
 "00000000000000000000010010010110", -- 1173 FREE #<CONS 0 1174>
 "00000000000000000000010010010111", -- 1174 FREE #<CONS 0 1175>
 "00000000000000000000010010011000", -- 1175 FREE #<CONS 0 1176>
 "00000000000000000000010010011001", -- 1176 FREE #<CONS 0 1177>
 "00000000000000000000010010011010", -- 1177 FREE #<CONS 0 1178>
 "00000000000000000000010010011011", -- 1178 FREE #<CONS 0 1179>
 "00000000000000000000010010011100", -- 1179 FREE #<CONS 0 1180>
 "00000000000000000000010010011101", -- 1180 FREE #<CONS 0 1181>
 "00000000000000000000010010011110", -- 1181 FREE #<CONS 0 1182>
 "00000000000000000000010010011111", -- 1182 FREE #<CONS 0 1183>
 "00000000000000000000010010100000", -- 1183 FREE #<CONS 0 1184>
 "00000000000000000000010010100001", -- 1184 FREE #<CONS 0 1185>
 "00000000000000000000010010100010", -- 1185 FREE #<CONS 0 1186>
 "00000000000000000000010010100011", -- 1186 FREE #<CONS 0 1187>
 "00000000000000000000010010100100", -- 1187 FREE #<CONS 0 1188>
 "00000000000000000000010010100101", -- 1188 FREE #<CONS 0 1189>
 "00000000000000000000010010100110", -- 1189 FREE #<CONS 0 1190>
 "00000000000000000000010010100111", -- 1190 FREE #<CONS 0 1191>
 "00000000000000000000010010101000", -- 1191 FREE #<CONS 0 1192>
 "00000000000000000000010010101001", -- 1192 FREE #<CONS 0 1193>
 "00000000000000000000010010101010", -- 1193 FREE #<CONS 0 1194>
 "00000000000000000000010010101011", -- 1194 FREE #<CONS 0 1195>
 "00000000000000000000010010101100", -- 1195 FREE #<CONS 0 1196>
 "00000000000000000000010010101101", -- 1196 FREE #<CONS 0 1197>
 "00000000000000000000010010101110", -- 1197 FREE #<CONS 0 1198>
 "00000000000000000000010010101111", -- 1198 FREE #<CONS 0 1199>
 "00000000000000000000010010110000", -- 1199 FREE #<CONS 0 1200>
 "00000000000000000000010010110001", -- 1200 FREE #<CONS 0 1201>
 "00000000000000000000010010110010", -- 1201 FREE #<CONS 0 1202>
 "00000000000000000000010010110011", -- 1202 FREE #<CONS 0 1203>
 "00000000000000000000010010110100", -- 1203 FREE #<CONS 0 1204>
 "00000000000000000000010010110101", -- 1204 FREE #<CONS 0 1205>
 "00000000000000000000010010110110", -- 1205 FREE #<CONS 0 1206>
 "00000000000000000000010010110111", -- 1206 FREE #<CONS 0 1207>
 "00000000000000000000010010111000", -- 1207 FREE #<CONS 0 1208>
 "00000000000000000000010010111001", -- 1208 FREE #<CONS 0 1209>
 "00000000000000000000010010111010", -- 1209 FREE #<CONS 0 1210>
 "00000000000000000000010010111011", -- 1210 FREE #<CONS 0 1211>
 "00000000000000000000010010111100", -- 1211 FREE #<CONS 0 1212>
 "00000000000000000000010010111101", -- 1212 FREE #<CONS 0 1213>
 "00000000000000000000010010111110", -- 1213 FREE #<CONS 0 1214>
 "00000000000000000000010010111111", -- 1214 FREE #<CONS 0 1215>
 "00000000000000000000010011000000", -- 1215 FREE #<CONS 0 1216>
 "00000000000000000000010011000001", -- 1216 FREE #<CONS 0 1217>
 "00000000000000000000010011000010", -- 1217 FREE #<CONS 0 1218>
 "00000000000000000000010011000011", -- 1218 FREE #<CONS 0 1219>
 "00000000000000000000010011000100", -- 1219 FREE #<CONS 0 1220>
 "00000000000000000000010011000101", -- 1220 FREE #<CONS 0 1221>
 "00000000000000000000010011000110", -- 1221 FREE #<CONS 0 1222>
 "00000000000000000000010011000111", -- 1222 FREE #<CONS 0 1223>
 "00000000000000000000010011001000", -- 1223 FREE #<CONS 0 1224>
 "00000000000000000000010011001001", -- 1224 FREE #<CONS 0 1225>
 "00000000000000000000010011001010", -- 1225 FREE #<CONS 0 1226>
 "00000000000000000000010011001011", -- 1226 FREE #<CONS 0 1227>
 "00000000000000000000010011001100", -- 1227 FREE #<CONS 0 1228>
 "00000000000000000000010011001101", -- 1228 FREE #<CONS 0 1229>
 "00000000000000000000010011001110", -- 1229 FREE #<CONS 0 1230>
 "00000000000000000000010011001111", -- 1230 FREE #<CONS 0 1231>
 "00000000000000000000010011010000", -- 1231 FREE #<CONS 0 1232>
 "00000000000000000000010011010001", -- 1232 FREE #<CONS 0 1233>
 "00000000000000000000010011010010", -- 1233 FREE #<CONS 0 1234>
 "00000000000000000000010011010011", -- 1234 FREE #<CONS 0 1235>
 "00000000000000000000010011010100", -- 1235 FREE #<CONS 0 1236>
 "00000000000000000000010011010101", -- 1236 FREE #<CONS 0 1237>
 "00000000000000000000010011010110", -- 1237 FREE #<CONS 0 1238>
 "00000000000000000000010011010111", -- 1238 FREE #<CONS 0 1239>
 "00000000000000000000010011011000", -- 1239 FREE #<CONS 0 1240>
 "00000000000000000000010011011001", -- 1240 FREE #<CONS 0 1241>
 "00000000000000000000010011011010", -- 1241 FREE #<CONS 0 1242>
 "00000000000000000000010011011011", -- 1242 FREE #<CONS 0 1243>
 "00000000000000000000010011011100", -- 1243 FREE #<CONS 0 1244>
 "00000000000000000000010011011101", -- 1244 FREE #<CONS 0 1245>
 "00000000000000000000010011011110", -- 1245 FREE #<CONS 0 1246>
 "00000000000000000000010011011111", -- 1246 FREE #<CONS 0 1247>
 "00000000000000000000010011100000", -- 1247 FREE #<CONS 0 1248>
 "00000000000000000000010011100001", -- 1248 FREE #<CONS 0 1249>
 "00000000000000000000010011100010", -- 1249 FREE #<CONS 0 1250>
 "00000000000000000000010011100011", -- 1250 FREE #<CONS 0 1251>
 "00000000000000000000010011100100", -- 1251 FREE #<CONS 0 1252>
 "00000000000000000000010011100101", -- 1252 FREE #<CONS 0 1253>
 "00000000000000000000010011100110", -- 1253 FREE #<CONS 0 1254>
 "00000000000000000000010011100111", -- 1254 FREE #<CONS 0 1255>
 "00000000000000000000010011101000", -- 1255 FREE #<CONS 0 1256>
 "00000000000000000000010011101001", -- 1256 FREE #<CONS 0 1257>
 "00000000000000000000010011101010", -- 1257 FREE #<CONS 0 1258>
 "00000000000000000000010011101011", -- 1258 FREE #<CONS 0 1259>
 "00000000000000000000010011101100", -- 1259 FREE #<CONS 0 1260>
 "00000000000000000000010011101101", -- 1260 FREE #<CONS 0 1261>
 "00000000000000000000010011101110", -- 1261 FREE #<CONS 0 1262>
 "00000000000000000000010011101111", -- 1262 FREE #<CONS 0 1263>
 "00000000000000000000010011110000", -- 1263 FREE #<CONS 0 1264>
 "00000000000000000000010011110001", -- 1264 FREE #<CONS 0 1265>
 "00000000000000000000010011110010", -- 1265 FREE #<CONS 0 1266>
 "00000000000000000000010011110011", -- 1266 FREE #<CONS 0 1267>
 "00000000000000000000010011110100", -- 1267 FREE #<CONS 0 1268>
 "00000000000000000000010011110101", -- 1268 FREE #<CONS 0 1269>
 "00000000000000000000010011110110", -- 1269 FREE #<CONS 0 1270>
 "00000000000000000000010011110111", -- 1270 FREE #<CONS 0 1271>
 "00000000000000000000010011111000", -- 1271 FREE #<CONS 0 1272>
 "00000000000000000000010011111001", -- 1272 FREE #<CONS 0 1273>
 "00000000000000000000010011111010", -- 1273 FREE #<CONS 0 1274>
 "00000000000000000000010011111011", -- 1274 FREE #<CONS 0 1275>
 "00000000000000000000010011111100", -- 1275 FREE #<CONS 0 1276>
 "00000000000000000000010011111101", -- 1276 FREE #<CONS 0 1277>
 "00000000000000000000010011111110", -- 1277 FREE #<CONS 0 1278>
 "00000000000000000000010011111111", -- 1278 FREE #<CONS 0 1279>
 "00000000000000000000010100000000", -- 1279 FREE #<CONS 0 1280>
 "00000000000000000000010100000001", -- 1280 FREE #<CONS 0 1281>
 "00000000000000000000010100000010", -- 1281 FREE #<CONS 0 1282>
 "00000000000000000000010100000011", -- 1282 FREE #<CONS 0 1283>
 "00000000000000000000010100000100", -- 1283 FREE #<CONS 0 1284>
 "00000000000000000000010100000101", -- 1284 FREE #<CONS 0 1285>
 "00000000000000000000010100000110", -- 1285 FREE #<CONS 0 1286>
 "00000000000000000000010100000111", -- 1286 FREE #<CONS 0 1287>
 "00000000000000000000010100001000", -- 1287 FREE #<CONS 0 1288>
 "00000000000000000000010100001001", -- 1288 FREE #<CONS 0 1289>
 "00000000000000000000010100001010", -- 1289 FREE #<CONS 0 1290>
 "00000000000000000000010100001011", -- 1290 FREE #<CONS 0 1291>
 "00000000000000000000010100001100", -- 1291 FREE #<CONS 0 1292>
 "00000000000000000000010100001101", -- 1292 FREE #<CONS 0 1293>
 "00000000000000000000010100001110", -- 1293 FREE #<CONS 0 1294>
 "00000000000000000000010100001111", -- 1294 FREE #<CONS 0 1295>
 "00000000000000000000010100010000", -- 1295 FREE #<CONS 0 1296>
 "00000000000000000000010100010001", -- 1296 FREE #<CONS 0 1297>
 "00000000000000000000010100010010", -- 1297 FREE #<CONS 0 1298>
 "00000000000000000000010100010011", -- 1298 FREE #<CONS 0 1299>
 "00000000000000000000010100010100", -- 1299 FREE #<CONS 0 1300>
 "00000000000000000000010100010101", -- 1300 FREE #<CONS 0 1301>
 "00000000000000000000010100010110", -- 1301 FREE #<CONS 0 1302>
 "00000000000000000000010100010111", -- 1302 FREE #<CONS 0 1303>
 "00000000000000000000010100011000", -- 1303 FREE #<CONS 0 1304>
 "00000000000000000000010100011001", -- 1304 FREE #<CONS 0 1305>
 "00000000000000000000010100011010", -- 1305 FREE #<CONS 0 1306>
 "00000000000000000000010100011011", -- 1306 FREE #<CONS 0 1307>
 "00000000000000000000010100011100", -- 1307 FREE #<CONS 0 1308>
 "00000000000000000000010100011101", -- 1308 FREE #<CONS 0 1309>
 "00000000000000000000010100011110", -- 1309 FREE #<CONS 0 1310>
 "00000000000000000000010100011111", -- 1310 FREE #<CONS 0 1311>
 "00000000000000000000010100100000", -- 1311 FREE #<CONS 0 1312>
 "00000000000000000000010100100001", -- 1312 FREE #<CONS 0 1313>
 "00000000000000000000010100100010", -- 1313 FREE #<CONS 0 1314>
 "00000000000000000000010100100011", -- 1314 FREE #<CONS 0 1315>
 "00000000000000000000010100100100", -- 1315 FREE #<CONS 0 1316>
 "00000000000000000000010100100101", -- 1316 FREE #<CONS 0 1317>
 "00000000000000000000010100100110", -- 1317 FREE #<CONS 0 1318>
 "00000000000000000000010100100111", -- 1318 FREE #<CONS 0 1319>
 "00000000000000000000010100101000", -- 1319 FREE #<CONS 0 1320>
 "00000000000000000000010100101001", -- 1320 FREE #<CONS 0 1321>
 "00000000000000000000010100101010", -- 1321 FREE #<CONS 0 1322>
 "00000000000000000000010100101011", -- 1322 FREE #<CONS 0 1323>
 "00000000000000000000010100101100", -- 1323 FREE #<CONS 0 1324>
 "00000000000000000000010100101101", -- 1324 FREE #<CONS 0 1325>
 "00000000000000000000010100101110", -- 1325 FREE #<CONS 0 1326>
 "00000000000000000000010100101111", -- 1326 FREE #<CONS 0 1327>
 "00000000000000000000010100110000", -- 1327 FREE #<CONS 0 1328>
 "00000000000000000000010100110001", -- 1328 FREE #<CONS 0 1329>
 "00000000000000000000010100110010", -- 1329 FREE #<CONS 0 1330>
 "00000000000000000000010100110011", -- 1330 FREE #<CONS 0 1331>
 "00000000000000000000010100110100", -- 1331 FREE #<CONS 0 1332>
 "00000000000000000000010100110101", -- 1332 FREE #<CONS 0 1333>
 "00000000000000000000010100110110", -- 1333 FREE #<CONS 0 1334>
 "00000000000000000000010100110111", -- 1334 FREE #<CONS 0 1335>
 "00000000000000000000010100111000", -- 1335 FREE #<CONS 0 1336>
 "00000000000000000000010100111001", -- 1336 FREE #<CONS 0 1337>
 "00000000000000000000010100111010", -- 1337 FREE #<CONS 0 1338>
 "00000000000000000000010100111011", -- 1338 FREE #<CONS 0 1339>
 "00000000000000000000010100111100", -- 1339 FREE #<CONS 0 1340>
 "00000000000000000000010100111101", -- 1340 FREE #<CONS 0 1341>
 "00000000000000000000010100111110", -- 1341 FREE #<CONS 0 1342>
 "00000000000000000000010100111111", -- 1342 FREE #<CONS 0 1343>
 "00000000000000000000010101000000", -- 1343 FREE #<CONS 0 1344>
 "00000000000000000000010101000001", -- 1344 FREE #<CONS 0 1345>
 "00000000000000000000010101000010", -- 1345 FREE #<CONS 0 1346>
 "00000000000000000000010101000011", -- 1346 FREE #<CONS 0 1347>
 "00000000000000000000010101000100", -- 1347 FREE #<CONS 0 1348>
 "00000000000000000000010101000101", -- 1348 FREE #<CONS 0 1349>
 "00000000000000000000010101000110", -- 1349 FREE #<CONS 0 1350>
 "00000000000000000000010101000111", -- 1350 FREE #<CONS 0 1351>
 "00000000000000000000010101001000", -- 1351 FREE #<CONS 0 1352>
 "00000000000000000000010101001001", -- 1352 FREE #<CONS 0 1353>
 "00000000000000000000010101001010", -- 1353 FREE #<CONS 0 1354>
 "00000000000000000000010101001011", -- 1354 FREE #<CONS 0 1355>
 "00000000000000000000010101001100", -- 1355 FREE #<CONS 0 1356>
 "00000000000000000000010101001101", -- 1356 FREE #<CONS 0 1357>
 "00000000000000000000010101001110", -- 1357 FREE #<CONS 0 1358>
 "00000000000000000000010101001111", -- 1358 FREE #<CONS 0 1359>
 "00000000000000000000010101010000", -- 1359 FREE #<CONS 0 1360>
 "00000000000000000000010101010001", -- 1360 FREE #<CONS 0 1361>
 "00000000000000000000010101010010", -- 1361 FREE #<CONS 0 1362>
 "00000000000000000000010101010011", -- 1362 FREE #<CONS 0 1363>
 "00000000000000000000010101010100", -- 1363 FREE #<CONS 0 1364>
 "00000000000000000000010101010101", -- 1364 FREE #<CONS 0 1365>
 "00000000000000000000010101010110", -- 1365 FREE #<CONS 0 1366>
 "00000000000000000000010101010111", -- 1366 FREE #<CONS 0 1367>
 "00000000000000000000010101011000", -- 1367 FREE #<CONS 0 1368>
 "00000000000000000000010101011001", -- 1368 FREE #<CONS 0 1369>
 "00000000000000000000010101011010", -- 1369 FREE #<CONS 0 1370>
 "00000000000000000000010101011011", -- 1370 FREE #<CONS 0 1371>
 "00000000000000000000010101011100", -- 1371 FREE #<CONS 0 1372>
 "00000000000000000000010101011101", -- 1372 FREE #<CONS 0 1373>
 "00000000000000000000010101011110", -- 1373 FREE #<CONS 0 1374>
 "00000000000000000000010101011111", -- 1374 FREE #<CONS 0 1375>
 "00000000000000000000010101100000", -- 1375 FREE #<CONS 0 1376>
 "00000000000000000000010101100001", -- 1376 FREE #<CONS 0 1377>
 "00000000000000000000010101100010", -- 1377 FREE #<CONS 0 1378>
 "00000000000000000000010101100011", -- 1378 FREE #<CONS 0 1379>
 "00000000000000000000010101100100", -- 1379 FREE #<CONS 0 1380>
 "00000000000000000000010101100101", -- 1380 FREE #<CONS 0 1381>
 "00000000000000000000010101100110", -- 1381 FREE #<CONS 0 1382>
 "00000000000000000000010101100111", -- 1382 FREE #<CONS 0 1383>
 "00000000000000000000010101101000", -- 1383 FREE #<CONS 0 1384>
 "00000000000000000000010101101001", -- 1384 FREE #<CONS 0 1385>
 "00000000000000000000010101101010", -- 1385 FREE #<CONS 0 1386>
 "00000000000000000000010101101011", -- 1386 FREE #<CONS 0 1387>
 "00000000000000000000010101101100", -- 1387 FREE #<CONS 0 1388>
 "00000000000000000000010101101101", -- 1388 FREE #<CONS 0 1389>
 "00000000000000000000010101101110", -- 1389 FREE #<CONS 0 1390>
 "00000000000000000000010101101111", -- 1390 FREE #<CONS 0 1391>
 "00000000000000000000010101110000", -- 1391 FREE #<CONS 0 1392>
 "00000000000000000000010101110001", -- 1392 FREE #<CONS 0 1393>
 "00000000000000000000010101110010", -- 1393 FREE #<CONS 0 1394>
 "00000000000000000000010101110011", -- 1394 FREE #<CONS 0 1395>
 "00000000000000000000010101110100", -- 1395 FREE #<CONS 0 1396>
 "00000000000000000000010101110101", -- 1396 FREE #<CONS 0 1397>
 "00000000000000000000010101110110", -- 1397 FREE #<CONS 0 1398>
 "00000000000000000000010101110111", -- 1398 FREE #<CONS 0 1399>
 "00000000000000000000010101111000", -- 1399 FREE #<CONS 0 1400>
 "00000000000000000000010101111001", -- 1400 FREE #<CONS 0 1401>
 "00000000000000000000010101111010", -- 1401 FREE #<CONS 0 1402>
 "00000000000000000000010101111011", -- 1402 FREE #<CONS 0 1403>
 "00000000000000000000010101111100", -- 1403 FREE #<CONS 0 1404>
 "00000000000000000000010101111101", -- 1404 FREE #<CONS 0 1405>
 "00000000000000000000010101111110", -- 1405 FREE #<CONS 0 1406>
 "00000000000000000000010101111111", -- 1406 FREE #<CONS 0 1407>
 "00000000000000000000010110000000", -- 1407 FREE #<CONS 0 1408>
 "00000000000000000000010110000001", -- 1408 FREE #<CONS 0 1409>
 "00000000000000000000010110000010", -- 1409 FREE #<CONS 0 1410>
 "00000000000000000000010110000011", -- 1410 FREE #<CONS 0 1411>
 "00000000000000000000010110000100", -- 1411 FREE #<CONS 0 1412>
 "00000000000000000000010110000101", -- 1412 FREE #<CONS 0 1413>
 "00000000000000000000010110000110", -- 1413 FREE #<CONS 0 1414>
 "00000000000000000000010110000111", -- 1414 FREE #<CONS 0 1415>
 "00000000000000000000010110001000", -- 1415 FREE #<CONS 0 1416>
 "00000000000000000000010110001001", -- 1416 FREE #<CONS 0 1417>
 "00000000000000000000010110001010", -- 1417 FREE #<CONS 0 1418>
 "00000000000000000000010110001011", -- 1418 FREE #<CONS 0 1419>
 "00000000000000000000010110001100", -- 1419 FREE #<CONS 0 1420>
 "00000000000000000000010110001101", -- 1420 FREE #<CONS 0 1421>
 "00000000000000000000010110001110", -- 1421 FREE #<CONS 0 1422>
 "00000000000000000000010110001111", -- 1422 FREE #<CONS 0 1423>
 "00000000000000000000010110010000", -- 1423 FREE #<CONS 0 1424>
 "00000000000000000000010110010001", -- 1424 FREE #<CONS 0 1425>
 "00000000000000000000010110010010", -- 1425 FREE #<CONS 0 1426>
 "00000000000000000000010110010011", -- 1426 FREE #<CONS 0 1427>
 "00000000000000000000010110010100", -- 1427 FREE #<CONS 0 1428>
 "00000000000000000000010110010101", -- 1428 FREE #<CONS 0 1429>
 "00000000000000000000010110010110", -- 1429 FREE #<CONS 0 1430>
 "00000000000000000000010110010111", -- 1430 FREE #<CONS 0 1431>
 "00000000000000000000010110011000", -- 1431 FREE #<CONS 0 1432>
 "00000000000000000000010110011001", -- 1432 FREE #<CONS 0 1433>
 "00000000000000000000010110011010", -- 1433 FREE #<CONS 0 1434>
 "00000000000000000000010110011011", -- 1434 FREE #<CONS 0 1435>
 "00000000000000000000010110011100", -- 1435 FREE #<CONS 0 1436>
 "00000000000000000000010110011101", -- 1436 FREE #<CONS 0 1437>
 "00000000000000000000010110011110", -- 1437 FREE #<CONS 0 1438>
 "00000000000000000000010110011111", -- 1438 FREE #<CONS 0 1439>
 "00000000000000000000010110100000", -- 1439 FREE #<CONS 0 1440>
 "00000000000000000000010110100001", -- 1440 FREE #<CONS 0 1441>
 "00000000000000000000010110100010", -- 1441 FREE #<CONS 0 1442>
 "00000000000000000000010110100011", -- 1442 FREE #<CONS 0 1443>
 "00000000000000000000010110100100", -- 1443 FREE #<CONS 0 1444>
 "00000000000000000000010110100101", -- 1444 FREE #<CONS 0 1445>
 "00000000000000000000010110100110", -- 1445 FREE #<CONS 0 1446>
 "00000000000000000000010110100111", -- 1446 FREE #<CONS 0 1447>
 "00000000000000000000010110101000", -- 1447 FREE #<CONS 0 1448>
 "00000000000000000000010110101001", -- 1448 FREE #<CONS 0 1449>
 "00000000000000000000010110101010", -- 1449 FREE #<CONS 0 1450>
 "00000000000000000000010110101011", -- 1450 FREE #<CONS 0 1451>
 "00000000000000000000010110101100", -- 1451 FREE #<CONS 0 1452>
 "00000000000000000000010110101101", -- 1452 FREE #<CONS 0 1453>
 "00000000000000000000010110101110", -- 1453 FREE #<CONS 0 1454>
 "00000000000000000000010110101111", -- 1454 FREE #<CONS 0 1455>
 "00000000000000000000010110110000", -- 1455 FREE #<CONS 0 1456>
 "00000000000000000000010110110001", -- 1456 FREE #<CONS 0 1457>
 "00000000000000000000010110110010", -- 1457 FREE #<CONS 0 1458>
 "00000000000000000000010110110011", -- 1458 FREE #<CONS 0 1459>
 "00000000000000000000010110110100", -- 1459 FREE #<CONS 0 1460>
 "00000000000000000000010110110101", -- 1460 FREE #<CONS 0 1461>
 "00000000000000000000010110110110", -- 1461 FREE #<CONS 0 1462>
 "00000000000000000000010110110111", -- 1462 FREE #<CONS 0 1463>
 "00000000000000000000010110111000", -- 1463 FREE #<CONS 0 1464>
 "00000000000000000000010110111001", -- 1464 FREE #<CONS 0 1465>
 "00000000000000000000010110111010", -- 1465 FREE #<CONS 0 1466>
 "00000000000000000000010110111011", -- 1466 FREE #<CONS 0 1467>
 "00000000000000000000010110111100", -- 1467 FREE #<CONS 0 1468>
 "00000000000000000000010110111101", -- 1468 FREE #<CONS 0 1469>
 "00000000000000000000010110111110", -- 1469 FREE #<CONS 0 1470>
 "00000000000000000000010110111111", -- 1470 FREE #<CONS 0 1471>
 "00000000000000000000010111000000", -- 1471 FREE #<CONS 0 1472>
 "00000000000000000000010111000001", -- 1472 FREE #<CONS 0 1473>
 "00000000000000000000010111000010", -- 1473 FREE #<CONS 0 1474>
 "00000000000000000000010111000011", -- 1474 FREE #<CONS 0 1475>
 "00000000000000000000010111000100", -- 1475 FREE #<CONS 0 1476>
 "00000000000000000000010111000101", -- 1476 FREE #<CONS 0 1477>
 "00000000000000000000010111000110", -- 1477 FREE #<CONS 0 1478>
 "00000000000000000000010111000111", -- 1478 FREE #<CONS 0 1479>
 "00000000000000000000010111001000", -- 1479 FREE #<CONS 0 1480>
 "00000000000000000000010111001001", -- 1480 FREE #<CONS 0 1481>
 "00000000000000000000010111001010", -- 1481 FREE #<CONS 0 1482>
 "00000000000000000000010111001011", -- 1482 FREE #<CONS 0 1483>
 "00000000000000000000010111001100", -- 1483 FREE #<CONS 0 1484>
 "00000000000000000000010111001101", -- 1484 FREE #<CONS 0 1485>
 "00000000000000000000010111001110", -- 1485 FREE #<CONS 0 1486>
 "00000000000000000000010111001111", -- 1486 FREE #<CONS 0 1487>
 "00000000000000000000010111010000", -- 1487 FREE #<CONS 0 1488>
 "00000000000000000000010111010001", -- 1488 FREE #<CONS 0 1489>
 "00000000000000000000010111010010", -- 1489 FREE #<CONS 0 1490>
 "00000000000000000000010111010011", -- 1490 FREE #<CONS 0 1491>
 "00000000000000000000010111010100", -- 1491 FREE #<CONS 0 1492>
 "00000000000000000000010111010101", -- 1492 FREE #<CONS 0 1493>
 "00000000000000000000010111010110", -- 1493 FREE #<CONS 0 1494>
 "00000000000000000000010111010111", -- 1494 FREE #<CONS 0 1495>
 "00000000000000000000010111011000", -- 1495 FREE #<CONS 0 1496>
 "00000000000000000000010111011001", -- 1496 FREE #<CONS 0 1497>
 "00000000000000000000010111011010", -- 1497 FREE #<CONS 0 1498>
 "00000000000000000000010111011011", -- 1498 FREE #<CONS 0 1499>
 "00000000000000000000010111011100", -- 1499 FREE #<CONS 0 1500>
 "00000000000000000000010111011101", -- 1500 FREE #<CONS 0 1501>
 "00000000000000000000010111011110", -- 1501 FREE #<CONS 0 1502>
 "00000000000000000000010111011111", -- 1502 FREE #<CONS 0 1503>
 "00000000000000000000010111100000", -- 1503 FREE #<CONS 0 1504>
 "00000000000000000000010111100001", -- 1504 FREE #<CONS 0 1505>
 "00000000000000000000010111100010", -- 1505 FREE #<CONS 0 1506>
 "00000000000000000000010111100011", -- 1506 FREE #<CONS 0 1507>
 "00000000000000000000010111100100", -- 1507 FREE #<CONS 0 1508>
 "00000000000000000000010111100101", -- 1508 FREE #<CONS 0 1509>
 "00000000000000000000010111100110", -- 1509 FREE #<CONS 0 1510>
 "00000000000000000000010111100111", -- 1510 FREE #<CONS 0 1511>
 "00000000000000000000010111101000", -- 1511 FREE #<CONS 0 1512>
 "00000000000000000000010111101001", -- 1512 FREE #<CONS 0 1513>
 "00000000000000000000010111101010", -- 1513 FREE #<CONS 0 1514>
 "00000000000000000000010111101011", -- 1514 FREE #<CONS 0 1515>
 "00000000000000000000010111101100", -- 1515 FREE #<CONS 0 1516>
 "00000000000000000000010111101101", -- 1516 FREE #<CONS 0 1517>
 "00000000000000000000010111101110", -- 1517 FREE #<CONS 0 1518>
 "00000000000000000000010111101111", -- 1518 FREE #<CONS 0 1519>
 "00000000000000000000010111110000", -- 1519 FREE #<CONS 0 1520>
 "00000000000000000000010111110001", -- 1520 FREE #<CONS 0 1521>
 "00000000000000000000010111110010", -- 1521 FREE #<CONS 0 1522>
 "00000000000000000000010111110011", -- 1522 FREE #<CONS 0 1523>
 "00000000000000000000010111110100", -- 1523 FREE #<CONS 0 1524>
 "00000000000000000000010111110101", -- 1524 FREE #<CONS 0 1525>
 "00000000000000000000010111110110", -- 1525 FREE #<CONS 0 1526>
 "00000000000000000000010111110111", -- 1526 FREE #<CONS 0 1527>
 "00000000000000000000010111111000", -- 1527 FREE #<CONS 0 1528>
 "00000000000000000000010111111001", -- 1528 FREE #<CONS 0 1529>
 "00000000000000000000010111111010", -- 1529 FREE #<CONS 0 1530>
 "00000000000000000000010111111011", -- 1530 FREE #<CONS 0 1531>
 "00000000000000000000010111111100", -- 1531 FREE #<CONS 0 1532>
 "00000000000000000000010111111101", -- 1532 FREE #<CONS 0 1533>
 "00000000000000000000010111111110", -- 1533 FREE #<CONS 0 1534>
 "00000000000000000000010111111111", -- 1534 FREE #<CONS 0 1535>
 "00000000000000000000011000000000", -- 1535 FREE #<CONS 0 1536>
 "00000000000000000000011000000001", -- 1536 FREE #<CONS 0 1537>
 "00000000000000000000011000000010", -- 1537 FREE #<CONS 0 1538>
 "00000000000000000000011000000011", -- 1538 FREE #<CONS 0 1539>
 "00000000000000000000011000000100", -- 1539 FREE #<CONS 0 1540>
 "00000000000000000000011000000101", -- 1540 FREE #<CONS 0 1541>
 "00000000000000000000011000000110", -- 1541 FREE #<CONS 0 1542>
 "00000000000000000000011000000111", -- 1542 FREE #<CONS 0 1543>
 "00000000000000000000011000001000", -- 1543 FREE #<CONS 0 1544>
 "00000000000000000000011000001001", -- 1544 FREE #<CONS 0 1545>
 "00000000000000000000011000001010", -- 1545 FREE #<CONS 0 1546>
 "00000000000000000000011000001011", -- 1546 FREE #<CONS 0 1547>
 "00000000000000000000011000001100", -- 1547 FREE #<CONS 0 1548>
 "00000000000000000000011000001101", -- 1548 FREE #<CONS 0 1549>
 "00000000000000000000011000001110", -- 1549 FREE #<CONS 0 1550>
 "00000000000000000000011000001111", -- 1550 FREE #<CONS 0 1551>
 "00000000000000000000011000010000", -- 1551 FREE #<CONS 0 1552>
 "00000000000000000000011000010001", -- 1552 FREE #<CONS 0 1553>
 "00000000000000000000011000010010", -- 1553 FREE #<CONS 0 1554>
 "00000000000000000000011000010011", -- 1554 FREE #<CONS 0 1555>
 "00000000000000000000011000010100", -- 1555 FREE #<CONS 0 1556>
 "00000000000000000000011000010101", -- 1556 FREE #<CONS 0 1557>
 "00000000000000000000011000010110", -- 1557 FREE #<CONS 0 1558>
 "00000000000000000000011000010111", -- 1558 FREE #<CONS 0 1559>
 "00000000000000000000011000011000", -- 1559 FREE #<CONS 0 1560>
 "00000000000000000000011000011001", -- 1560 FREE #<CONS 0 1561>
 "00000000000000000000011000011010", -- 1561 FREE #<CONS 0 1562>
 "00000000000000000000011000011011", -- 1562 FREE #<CONS 0 1563>
 "00000000000000000000011000011100", -- 1563 FREE #<CONS 0 1564>
 "00000000000000000000011000011101", -- 1564 FREE #<CONS 0 1565>
 "00000000000000000000011000011110", -- 1565 FREE #<CONS 0 1566>
 "00000000000000000000011000011111", -- 1566 FREE #<CONS 0 1567>
 "00000000000000000000011000100000", -- 1567 FREE #<CONS 0 1568>
 "00000000000000000000011000100001", -- 1568 FREE #<CONS 0 1569>
 "00000000000000000000011000100010", -- 1569 FREE #<CONS 0 1570>
 "00000000000000000000011000100011", -- 1570 FREE #<CONS 0 1571>
 "00000000000000000000011000100100", -- 1571 FREE #<CONS 0 1572>
 "00000000000000000000011000100101", -- 1572 FREE #<CONS 0 1573>
 "00000000000000000000011000100110", -- 1573 FREE #<CONS 0 1574>
 "00000000000000000000011000100111", -- 1574 FREE #<CONS 0 1575>
 "00000000000000000000011000101000", -- 1575 FREE #<CONS 0 1576>
 "00000000000000000000011000101001", -- 1576 FREE #<CONS 0 1577>
 "00000000000000000000011000101010", -- 1577 FREE #<CONS 0 1578>
 "00000000000000000000011000101011", -- 1578 FREE #<CONS 0 1579>
 "00000000000000000000011000101100", -- 1579 FREE #<CONS 0 1580>
 "00000000000000000000011000101101", -- 1580 FREE #<CONS 0 1581>
 "00000000000000000000011000101110", -- 1581 FREE #<CONS 0 1582>
 "00000000000000000000011000101111", -- 1582 FREE #<CONS 0 1583>
 "00000000000000000000011000110000", -- 1583 FREE #<CONS 0 1584>
 "00000000000000000000011000110001", -- 1584 FREE #<CONS 0 1585>
 "00000000000000000000011000110010", -- 1585 FREE #<CONS 0 1586>
 "00000000000000000000011000110011", -- 1586 FREE #<CONS 0 1587>
 "00000000000000000000011000110100", -- 1587 FREE #<CONS 0 1588>
 "00000000000000000000011000110101", -- 1588 FREE #<CONS 0 1589>
 "00000000000000000000011000110110", -- 1589 FREE #<CONS 0 1590>
 "00000000000000000000011000110111", -- 1590 FREE #<CONS 0 1591>
 "00000000000000000000011000111000", -- 1591 FREE #<CONS 0 1592>
 "00000000000000000000011000111001", -- 1592 FREE #<CONS 0 1593>
 "00000000000000000000011000111010", -- 1593 FREE #<CONS 0 1594>
 "00000000000000000000011000111011", -- 1594 FREE #<CONS 0 1595>
 "00000000000000000000011000111100", -- 1595 FREE #<CONS 0 1596>
 "00000000000000000000011000111101", -- 1596 FREE #<CONS 0 1597>
 "00000000000000000000011000111110", -- 1597 FREE #<CONS 0 1598>
 "00000000000000000000011000111111", -- 1598 FREE #<CONS 0 1599>
 "00000000000000000000011001000000", -- 1599 FREE #<CONS 0 1600>
 "00000000000000000000011001000001", -- 1600 FREE #<CONS 0 1601>
 "00000000000000000000011001000010", -- 1601 FREE #<CONS 0 1602>
 "00000000000000000000011001000011", -- 1602 FREE #<CONS 0 1603>
 "00000000000000000000011001000100", -- 1603 FREE #<CONS 0 1604>
 "00000000000000000000011001000101", -- 1604 FREE #<CONS 0 1605>
 "00000000000000000000011001000110", -- 1605 FREE #<CONS 0 1606>
 "00000000000000000000011001000111", -- 1606 FREE #<CONS 0 1607>
 "00000000000000000000011001001000", -- 1607 FREE #<CONS 0 1608>
 "00000000000000000000011001001001", -- 1608 FREE #<CONS 0 1609>
 "00000000000000000000011001001010", -- 1609 FREE #<CONS 0 1610>
 "00000000000000000000011001001011", -- 1610 FREE #<CONS 0 1611>
 "00000000000000000000011001001100", -- 1611 FREE #<CONS 0 1612>
 "00000000000000000000011001001101", -- 1612 FREE #<CONS 0 1613>
 "00000000000000000000011001001110", -- 1613 FREE #<CONS 0 1614>
 "00000000000000000000011001001111", -- 1614 FREE #<CONS 0 1615>
 "00000000000000000000011001010000", -- 1615 FREE #<CONS 0 1616>
 "00000000000000000000011001010001", -- 1616 FREE #<CONS 0 1617>
 "00000000000000000000011001010010", -- 1617 FREE #<CONS 0 1618>
 "00000000000000000000011001010011", -- 1618 FREE #<CONS 0 1619>
 "00000000000000000000011001010100", -- 1619 FREE #<CONS 0 1620>
 "00000000000000000000011001010101", -- 1620 FREE #<CONS 0 1621>
 "00000000000000000000011001010110", -- 1621 FREE #<CONS 0 1622>
 "00000000000000000000011001010111", -- 1622 FREE #<CONS 0 1623>
 "00000000000000000000011001011000", -- 1623 FREE #<CONS 0 1624>
 "00000000000000000000011001011001", -- 1624 FREE #<CONS 0 1625>
 "00000000000000000000011001011010", -- 1625 FREE #<CONS 0 1626>
 "00000000000000000000011001011011", -- 1626 FREE #<CONS 0 1627>
 "00000000000000000000011001011100", -- 1627 FREE #<CONS 0 1628>
 "00000000000000000000011001011101", -- 1628 FREE #<CONS 0 1629>
 "00000000000000000000011001011110", -- 1629 FREE #<CONS 0 1630>
 "00000000000000000000011001011111", -- 1630 FREE #<CONS 0 1631>
 "00000000000000000000011001100000", -- 1631 FREE #<CONS 0 1632>
 "00000000000000000000011001100001", -- 1632 FREE #<CONS 0 1633>
 "00000000000000000000011001100010", -- 1633 FREE #<CONS 0 1634>
 "00000000000000000000011001100011", -- 1634 FREE #<CONS 0 1635>
 "00000000000000000000011001100100", -- 1635 FREE #<CONS 0 1636>
 "00000000000000000000011001100101", -- 1636 FREE #<CONS 0 1637>
 "00000000000000000000011001100110", -- 1637 FREE #<CONS 0 1638>
 "00000000000000000000011001100111", -- 1638 FREE #<CONS 0 1639>
 "00000000000000000000011001101000", -- 1639 FREE #<CONS 0 1640>
 "00000000000000000000011001101001", -- 1640 FREE #<CONS 0 1641>
 "00000000000000000000011001101010", -- 1641 FREE #<CONS 0 1642>
 "00000000000000000000011001101011", -- 1642 FREE #<CONS 0 1643>
 "00000000000000000000011001101100", -- 1643 FREE #<CONS 0 1644>
 "00000000000000000000011001101101", -- 1644 FREE #<CONS 0 1645>
 "00000000000000000000011001101110", -- 1645 FREE #<CONS 0 1646>
 "00000000000000000000011001101111", -- 1646 FREE #<CONS 0 1647>
 "00000000000000000000011001110000", -- 1647 FREE #<CONS 0 1648>
 "00000000000000000000011001110001", -- 1648 FREE #<CONS 0 1649>
 "00000000000000000000011001110010", -- 1649 FREE #<CONS 0 1650>
 "00000000000000000000011001110011", -- 1650 FREE #<CONS 0 1651>
 "00000000000000000000011001110100", -- 1651 FREE #<CONS 0 1652>
 "00000000000000000000011001110101", -- 1652 FREE #<CONS 0 1653>
 "00000000000000000000011001110110", -- 1653 FREE #<CONS 0 1654>
 "00000000000000000000011001110111", -- 1654 FREE #<CONS 0 1655>
 "00000000000000000000011001111000", -- 1655 FREE #<CONS 0 1656>
 "00000000000000000000011001111001", -- 1656 FREE #<CONS 0 1657>
 "00000000000000000000011001111010", -- 1657 FREE #<CONS 0 1658>
 "00000000000000000000011001111011", -- 1658 FREE #<CONS 0 1659>
 "00000000000000000000011001111100", -- 1659 FREE #<CONS 0 1660>
 "00000000000000000000011001111101", -- 1660 FREE #<CONS 0 1661>
 "00000000000000000000011001111110", -- 1661 FREE #<CONS 0 1662>
 "00000000000000000000011001111111", -- 1662 FREE #<CONS 0 1663>
 "00000000000000000000011010000000", -- 1663 FREE #<CONS 0 1664>
 "00000000000000000000011010000001", -- 1664 FREE #<CONS 0 1665>
 "00000000000000000000011010000010", -- 1665 FREE #<CONS 0 1666>
 "00000000000000000000011010000011", -- 1666 FREE #<CONS 0 1667>
 "00000000000000000000011010000100", -- 1667 FREE #<CONS 0 1668>
 "00000000000000000000011010000101", -- 1668 FREE #<CONS 0 1669>
 "00000000000000000000011010000110", -- 1669 FREE #<CONS 0 1670>
 "00000000000000000000011010000111", -- 1670 FREE #<CONS 0 1671>
 "00000000000000000000011010001000", -- 1671 FREE #<CONS 0 1672>
 "00000000000000000000011010001001", -- 1672 FREE #<CONS 0 1673>
 "00000000000000000000011010001010", -- 1673 FREE #<CONS 0 1674>
 "00000000000000000000011010001011", -- 1674 FREE #<CONS 0 1675>
 "00000000000000000000011010001100", -- 1675 FREE #<CONS 0 1676>
 "00000000000000000000011010001101", -- 1676 FREE #<CONS 0 1677>
 "00000000000000000000011010001110", -- 1677 FREE #<CONS 0 1678>
 "00000000000000000000011010001111", -- 1678 FREE #<CONS 0 1679>
 "00000000000000000000011010010000", -- 1679 FREE #<CONS 0 1680>
 "00000000000000000000011010010001", -- 1680 FREE #<CONS 0 1681>
 "00000000000000000000011010010010", -- 1681 FREE #<CONS 0 1682>
 "00000000000000000000011010010011", -- 1682 FREE #<CONS 0 1683>
 "00000000000000000000011010010100", -- 1683 FREE #<CONS 0 1684>
 "00000000000000000000011010010101", -- 1684 FREE #<CONS 0 1685>
 "00000000000000000000011010010110", -- 1685 FREE #<CONS 0 1686>
 "00000000000000000000011010010111", -- 1686 FREE #<CONS 0 1687>
 "00000000000000000000011010011000", -- 1687 FREE #<CONS 0 1688>
 "00000000000000000000011010011001", -- 1688 FREE #<CONS 0 1689>
 "00000000000000000000011010011010", -- 1689 FREE #<CONS 0 1690>
 "00000000000000000000011010011011", -- 1690 FREE #<CONS 0 1691>
 "00000000000000000000011010011100", -- 1691 FREE #<CONS 0 1692>
 "00000000000000000000011010011101", -- 1692 FREE #<CONS 0 1693>
 "00000000000000000000011010011110", -- 1693 FREE #<CONS 0 1694>
 "00000000000000000000011010011111", -- 1694 FREE #<CONS 0 1695>
 "00000000000000000000011010100000", -- 1695 FREE #<CONS 0 1696>
 "00000000000000000000011010100001", -- 1696 FREE #<CONS 0 1697>
 "00000000000000000000011010100010", -- 1697 FREE #<CONS 0 1698>
 "00000000000000000000011010100011", -- 1698 FREE #<CONS 0 1699>
 "00000000000000000000011010100100", -- 1699 FREE #<CONS 0 1700>
 "00000000000000000000011010100101", -- 1700 FREE #<CONS 0 1701>
 "00000000000000000000011010100110", -- 1701 FREE #<CONS 0 1702>
 "00000000000000000000011010100111", -- 1702 FREE #<CONS 0 1703>
 "00000000000000000000011010101000", -- 1703 FREE #<CONS 0 1704>
 "00000000000000000000011010101001", -- 1704 FREE #<CONS 0 1705>
 "00000000000000000000011010101010", -- 1705 FREE #<CONS 0 1706>
 "00000000000000000000011010101011", -- 1706 FREE #<CONS 0 1707>
 "00000000000000000000011010101100", -- 1707 FREE #<CONS 0 1708>
 "00000000000000000000011010101101", -- 1708 FREE #<CONS 0 1709>
 "00000000000000000000011010101110", -- 1709 FREE #<CONS 0 1710>
 "00000000000000000000011010101111", -- 1710 FREE #<CONS 0 1711>
 "00000000000000000000011010110000", -- 1711 FREE #<CONS 0 1712>
 "00000000000000000000011010110001", -- 1712 FREE #<CONS 0 1713>
 "00000000000000000000011010110010", -- 1713 FREE #<CONS 0 1714>
 "00000000000000000000011010110011", -- 1714 FREE #<CONS 0 1715>
 "00000000000000000000011010110100", -- 1715 FREE #<CONS 0 1716>
 "00000000000000000000011010110101", -- 1716 FREE #<CONS 0 1717>
 "00000000000000000000011010110110", -- 1717 FREE #<CONS 0 1718>
 "00000000000000000000011010110111", -- 1718 FREE #<CONS 0 1719>
 "00000000000000000000011010111000", -- 1719 FREE #<CONS 0 1720>
 "00000000000000000000011010111001", -- 1720 FREE #<CONS 0 1721>
 "00000000000000000000011010111010", -- 1721 FREE #<CONS 0 1722>
 "00000000000000000000011010111011", -- 1722 FREE #<CONS 0 1723>
 "00000000000000000000011010111100", -- 1723 FREE #<CONS 0 1724>
 "00000000000000000000011010111101", -- 1724 FREE #<CONS 0 1725>
 "00000000000000000000011010111110", -- 1725 FREE #<CONS 0 1726>
 "00000000000000000000011010111111", -- 1726 FREE #<CONS 0 1727>
 "00000000000000000000011011000000", -- 1727 FREE #<CONS 0 1728>
 "00000000000000000000011011000001", -- 1728 FREE #<CONS 0 1729>
 "00000000000000000000011011000010", -- 1729 FREE #<CONS 0 1730>
 "00000000000000000000011011000011", -- 1730 FREE #<CONS 0 1731>
 "00000000000000000000011011000100", -- 1731 FREE #<CONS 0 1732>
 "00000000000000000000011011000101", -- 1732 FREE #<CONS 0 1733>
 "00000000000000000000011011000110", -- 1733 FREE #<CONS 0 1734>
 "00000000000000000000011011000111", -- 1734 FREE #<CONS 0 1735>
 "00000000000000000000011011001000", -- 1735 FREE #<CONS 0 1736>
 "00000000000000000000011011001001", -- 1736 FREE #<CONS 0 1737>
 "00000000000000000000011011001010", -- 1737 FREE #<CONS 0 1738>
 "00000000000000000000011011001011", -- 1738 FREE #<CONS 0 1739>
 "00000000000000000000011011001100", -- 1739 FREE #<CONS 0 1740>
 "00000000000000000000011011001101", -- 1740 FREE #<CONS 0 1741>
 "00000000000000000000011011001110", -- 1741 FREE #<CONS 0 1742>
 "00000000000000000000011011001111", -- 1742 FREE #<CONS 0 1743>
 "00000000000000000000011011010000", -- 1743 FREE #<CONS 0 1744>
 "00000000000000000000011011010001", -- 1744 FREE #<CONS 0 1745>
 "00000000000000000000011011010010", -- 1745 FREE #<CONS 0 1746>
 "00000000000000000000011011010011", -- 1746 FREE #<CONS 0 1747>
 "00000000000000000000011011010100", -- 1747 FREE #<CONS 0 1748>
 "00000000000000000000011011010101", -- 1748 FREE #<CONS 0 1749>
 "00000000000000000000011011010110", -- 1749 FREE #<CONS 0 1750>
 "00000000000000000000011011010111", -- 1750 FREE #<CONS 0 1751>
 "00000000000000000000011011011000", -- 1751 FREE #<CONS 0 1752>
 "00000000000000000000011011011001", -- 1752 FREE #<CONS 0 1753>
 "00000000000000000000011011011010", -- 1753 FREE #<CONS 0 1754>
 "00000000000000000000011011011011", -- 1754 FREE #<CONS 0 1755>
 "00000000000000000000011011011100", -- 1755 FREE #<CONS 0 1756>
 "00000000000000000000011011011101", -- 1756 FREE #<CONS 0 1757>
 "00000000000000000000011011011110", -- 1757 FREE #<CONS 0 1758>
 "00000000000000000000011011011111", -- 1758 FREE #<CONS 0 1759>
 "00000000000000000000011011100000", -- 1759 FREE #<CONS 0 1760>
 "00000000000000000000011011100001", -- 1760 FREE #<CONS 0 1761>
 "00000000000000000000011011100010", -- 1761 FREE #<CONS 0 1762>
 "00000000000000000000011011100011", -- 1762 FREE #<CONS 0 1763>
 "00000000000000000000011011100100", -- 1763 FREE #<CONS 0 1764>
 "00000000000000000000011011100101", -- 1764 FREE #<CONS 0 1765>
 "00000000000000000000011011100110", -- 1765 FREE #<CONS 0 1766>
 "00000000000000000000011011100111", -- 1766 FREE #<CONS 0 1767>
 "00000000000000000000011011101000", -- 1767 FREE #<CONS 0 1768>
 "00000000000000000000011011101001", -- 1768 FREE #<CONS 0 1769>
 "00000000000000000000011011101010", -- 1769 FREE #<CONS 0 1770>
 "00000000000000000000011011101011", -- 1770 FREE #<CONS 0 1771>
 "00000000000000000000011011101100", -- 1771 FREE #<CONS 0 1772>
 "00000000000000000000011011101101", -- 1772 FREE #<CONS 0 1773>
 "00000000000000000000011011101110", -- 1773 FREE #<CONS 0 1774>
 "00000000000000000000011011101111", -- 1774 FREE #<CONS 0 1775>
 "00000000000000000000011011110000", -- 1775 FREE #<CONS 0 1776>
 "00000000000000000000011011110001", -- 1776 FREE #<CONS 0 1777>
 "00000000000000000000011011110010", -- 1777 FREE #<CONS 0 1778>
 "00000000000000000000011011110011", -- 1778 FREE #<CONS 0 1779>
 "00000000000000000000011011110100", -- 1779 FREE #<CONS 0 1780>
 "00000000000000000000011011110101", -- 1780 FREE #<CONS 0 1781>
 "00000000000000000000011011110110", -- 1781 FREE #<CONS 0 1782>
 "00000000000000000000011011110111", -- 1782 FREE #<CONS 0 1783>
 "00000000000000000000011011111000", -- 1783 FREE #<CONS 0 1784>
 "00000000000000000000011011111001", -- 1784 FREE #<CONS 0 1785>
 "00000000000000000000011011111010", -- 1785 FREE #<CONS 0 1786>
 "00000000000000000000011011111011", -- 1786 FREE #<CONS 0 1787>
 "00000000000000000000011011111100", -- 1787 FREE #<CONS 0 1788>
 "00000000000000000000011011111101", -- 1788 FREE #<CONS 0 1789>
 "00000000000000000000011011111110", -- 1789 FREE #<CONS 0 1790>
 "00000000000000000000011011111111", -- 1790 FREE #<CONS 0 1791>
 "00000000000000000000011100000000", -- 1791 FREE #<CONS 0 1792>
 "00000000000000000000011100000001", -- 1792 FREE #<CONS 0 1793>
 "00000000000000000000011100000010", -- 1793 FREE #<CONS 0 1794>
 "00000000000000000000011100000011", -- 1794 FREE #<CONS 0 1795>
 "00000000000000000000011100000100", -- 1795 FREE #<CONS 0 1796>
 "00000000000000000000011100000101", -- 1796 FREE #<CONS 0 1797>
 "00000000000000000000011100000110", -- 1797 FREE #<CONS 0 1798>
 "00000000000000000000011100000111", -- 1798 FREE #<CONS 0 1799>
 "00000000000000000000011100001000", -- 1799 FREE #<CONS 0 1800>
 "00000000000000000000011100001001", -- 1800 FREE #<CONS 0 1801>
 "00000000000000000000011100001010", -- 1801 FREE #<CONS 0 1802>
 "00000000000000000000011100001011", -- 1802 FREE #<CONS 0 1803>
 "00000000000000000000011100001100", -- 1803 FREE #<CONS 0 1804>
 "00000000000000000000011100001101", -- 1804 FREE #<CONS 0 1805>
 "00000000000000000000011100001110", -- 1805 FREE #<CONS 0 1806>
 "00000000000000000000011100001111", -- 1806 FREE #<CONS 0 1807>
 "00000000000000000000011100010000", -- 1807 FREE #<CONS 0 1808>
 "00000000000000000000011100010001", -- 1808 FREE #<CONS 0 1809>
 "00000000000000000000011100010010", -- 1809 FREE #<CONS 0 1810>
 "00000000000000000000011100010011", -- 1810 FREE #<CONS 0 1811>
 "00000000000000000000011100010100", -- 1811 FREE #<CONS 0 1812>
 "00000000000000000000011100010101", -- 1812 FREE #<CONS 0 1813>
 "00000000000000000000011100010110", -- 1813 FREE #<CONS 0 1814>
 "00000000000000000000011100010111", -- 1814 FREE #<CONS 0 1815>
 "00000000000000000000011100011000", -- 1815 FREE #<CONS 0 1816>
 "00000000000000000000011100011001", -- 1816 FREE #<CONS 0 1817>
 "00000000000000000000011100011010", -- 1817 FREE #<CONS 0 1818>
 "00000000000000000000011100011011", -- 1818 FREE #<CONS 0 1819>
 "00000000000000000000011100011100", -- 1819 FREE #<CONS 0 1820>
 "00000000000000000000011100011101", -- 1820 FREE #<CONS 0 1821>
 "00000000000000000000011100011110", -- 1821 FREE #<CONS 0 1822>
 "00000000000000000000011100011111", -- 1822 FREE #<CONS 0 1823>
 "00000000000000000000011100100000", -- 1823 FREE #<CONS 0 1824>
 "00000000000000000000011100100001", -- 1824 FREE #<CONS 0 1825>
 "00000000000000000000011100100010", -- 1825 FREE #<CONS 0 1826>
 "00000000000000000000011100100011", -- 1826 FREE #<CONS 0 1827>
 "00000000000000000000011100100100", -- 1827 FREE #<CONS 0 1828>
 "00000000000000000000011100100101", -- 1828 FREE #<CONS 0 1829>
 "00000000000000000000011100100110", -- 1829 FREE #<CONS 0 1830>
 "00000000000000000000011100100111", -- 1830 FREE #<CONS 0 1831>
 "00000000000000000000011100101000", -- 1831 FREE #<CONS 0 1832>
 "00000000000000000000011100101001", -- 1832 FREE #<CONS 0 1833>
 "00000000000000000000011100101010", -- 1833 FREE #<CONS 0 1834>
 "00000000000000000000011100101011", -- 1834 FREE #<CONS 0 1835>
 "00000000000000000000011100101100", -- 1835 FREE #<CONS 0 1836>
 "00000000000000000000011100101101", -- 1836 FREE #<CONS 0 1837>
 "00000000000000000000011100101110", -- 1837 FREE #<CONS 0 1838>
 "00000000000000000000011100101111", -- 1838 FREE #<CONS 0 1839>
 "00000000000000000000011100110000", -- 1839 FREE #<CONS 0 1840>
 "00000000000000000000011100110001", -- 1840 FREE #<CONS 0 1841>
 "00000000000000000000011100110010", -- 1841 FREE #<CONS 0 1842>
 "00000000000000000000011100110011", -- 1842 FREE #<CONS 0 1843>
 "00000000000000000000011100110100", -- 1843 FREE #<CONS 0 1844>
 "00000000000000000000011100110101", -- 1844 FREE #<CONS 0 1845>
 "00000000000000000000011100110110", -- 1845 FREE #<CONS 0 1846>
 "00000000000000000000011100110111", -- 1846 FREE #<CONS 0 1847>
 "00000000000000000000011100111000", -- 1847 FREE #<CONS 0 1848>
 "00000000000000000000011100111001", -- 1848 FREE #<CONS 0 1849>
 "00000000000000000000011100111010", -- 1849 FREE #<CONS 0 1850>
 "00000000000000000000011100111011", -- 1850 FREE #<CONS 0 1851>
 "00000000000000000000011100111100", -- 1851 FREE #<CONS 0 1852>
 "00000000000000000000011100111101", -- 1852 FREE #<CONS 0 1853>
 "00000000000000000000011100111110", -- 1853 FREE #<CONS 0 1854>
 "00000000000000000000011100111111", -- 1854 FREE #<CONS 0 1855>
 "00000000000000000000011101000000", -- 1855 FREE #<CONS 0 1856>
 "00000000000000000000011101000001", -- 1856 FREE #<CONS 0 1857>
 "00000000000000000000011101000010", -- 1857 FREE #<CONS 0 1858>
 "00000000000000000000011101000011", -- 1858 FREE #<CONS 0 1859>
 "00000000000000000000011101000100", -- 1859 FREE #<CONS 0 1860>
 "00000000000000000000011101000101", -- 1860 FREE #<CONS 0 1861>
 "00000000000000000000011101000110", -- 1861 FREE #<CONS 0 1862>
 "00000000000000000000011101000111", -- 1862 FREE #<CONS 0 1863>
 "00000000000000000000011101001000", -- 1863 FREE #<CONS 0 1864>
 "00000000000000000000011101001001", -- 1864 FREE #<CONS 0 1865>
 "00000000000000000000011101001010", -- 1865 FREE #<CONS 0 1866>
 "00000000000000000000011101001011", -- 1866 FREE #<CONS 0 1867>
 "00000000000000000000011101001100", -- 1867 FREE #<CONS 0 1868>
 "00000000000000000000011101001101", -- 1868 FREE #<CONS 0 1869>
 "00000000000000000000011101001110", -- 1869 FREE #<CONS 0 1870>
 "00000000000000000000011101001111", -- 1870 FREE #<CONS 0 1871>
 "00000000000000000000011101010000", -- 1871 FREE #<CONS 0 1872>
 "00000000000000000000011101010001", -- 1872 FREE #<CONS 0 1873>
 "00000000000000000000011101010010", -- 1873 FREE #<CONS 0 1874>
 "00000000000000000000011101010011", -- 1874 FREE #<CONS 0 1875>
 "00000000000000000000011101010100", -- 1875 FREE #<CONS 0 1876>
 "00000000000000000000011101010101", -- 1876 FREE #<CONS 0 1877>
 "00000000000000000000011101010110", -- 1877 FREE #<CONS 0 1878>
 "00000000000000000000011101010111", -- 1878 FREE #<CONS 0 1879>
 "00000000000000000000011101011000", -- 1879 FREE #<CONS 0 1880>
 "00000000000000000000011101011001", -- 1880 FREE #<CONS 0 1881>
 "00000000000000000000011101011010", -- 1881 FREE #<CONS 0 1882>
 "00000000000000000000011101011011", -- 1882 FREE #<CONS 0 1883>
 "00000000000000000000011101011100", -- 1883 FREE #<CONS 0 1884>
 "00000000000000000000011101011101", -- 1884 FREE #<CONS 0 1885>
 "00000000000000000000011101011110", -- 1885 FREE #<CONS 0 1886>
 "00000000000000000000011101011111", -- 1886 FREE #<CONS 0 1887>
 "00000000000000000000011101100000", -- 1887 FREE #<CONS 0 1888>
 "00000000000000000000011101100001", -- 1888 FREE #<CONS 0 1889>
 "00000000000000000000011101100010", -- 1889 FREE #<CONS 0 1890>
 "00000000000000000000011101100011", -- 1890 FREE #<CONS 0 1891>
 "00000000000000000000011101100100", -- 1891 FREE #<CONS 0 1892>
 "00000000000000000000011101100101", -- 1892 FREE #<CONS 0 1893>
 "00000000000000000000011101100110", -- 1893 FREE #<CONS 0 1894>
 "00000000000000000000011101100111", -- 1894 FREE #<CONS 0 1895>
 "00000000000000000000011101101000", -- 1895 FREE #<CONS 0 1896>
 "00000000000000000000011101101001", -- 1896 FREE #<CONS 0 1897>
 "00000000000000000000011101101010", -- 1897 FREE #<CONS 0 1898>
 "00000000000000000000011101101011", -- 1898 FREE #<CONS 0 1899>
 "00000000000000000000011101101100", -- 1899 FREE #<CONS 0 1900>
 "00000000000000000000011101101101", -- 1900 FREE #<CONS 0 1901>
 "00000000000000000000011101101110", -- 1901 FREE #<CONS 0 1902>
 "00000000000000000000011101101111", -- 1902 FREE #<CONS 0 1903>
 "00000000000000000000011101110000", -- 1903 FREE #<CONS 0 1904>
 "00000000000000000000011101110001", -- 1904 FREE #<CONS 0 1905>
 "00000000000000000000011101110010", -- 1905 FREE #<CONS 0 1906>
 "00000000000000000000011101110011", -- 1906 FREE #<CONS 0 1907>
 "00000000000000000000011101110100", -- 1907 FREE #<CONS 0 1908>
 "00000000000000000000011101110101", -- 1908 FREE #<CONS 0 1909>
 "00000000000000000000011101110110", -- 1909 FREE #<CONS 0 1910>
 "00000000000000000000011101110111", -- 1910 FREE #<CONS 0 1911>
 "00000000000000000000011101111000", -- 1911 FREE #<CONS 0 1912>
 "00000000000000000000011101111001", -- 1912 FREE #<CONS 0 1913>
 "00000000000000000000011101111010", -- 1913 FREE #<CONS 0 1914>
 "00000000000000000000011101111011", -- 1914 FREE #<CONS 0 1915>
 "00000000000000000000011101111100", -- 1915 FREE #<CONS 0 1916>
 "00000000000000000000011101111101", -- 1916 FREE #<CONS 0 1917>
 "00000000000000000000011101111110", -- 1917 FREE #<CONS 0 1918>
 "00000000000000000000011101111111", -- 1918 FREE #<CONS 0 1919>
 "00000000000000000000011110000000", -- 1919 FREE #<CONS 0 1920>
 "00000000000000000000011110000001", -- 1920 FREE #<CONS 0 1921>
 "00000000000000000000011110000010", -- 1921 FREE #<CONS 0 1922>
 "00000000000000000000011110000011", -- 1922 FREE #<CONS 0 1923>
 "00000000000000000000011110000100", -- 1923 FREE #<CONS 0 1924>
 "00000000000000000000011110000101", -- 1924 FREE #<CONS 0 1925>
 "00000000000000000000011110000110", -- 1925 FREE #<CONS 0 1926>
 "00000000000000000000011110000111", -- 1926 FREE #<CONS 0 1927>
 "00000000000000000000011110001000", -- 1927 FREE #<CONS 0 1928>
 "00000000000000000000011110001001", -- 1928 FREE #<CONS 0 1929>
 "00000000000000000000011110001010", -- 1929 FREE #<CONS 0 1930>
 "00000000000000000000011110001011", -- 1930 FREE #<CONS 0 1931>
 "00000000000000000000011110001100", -- 1931 FREE #<CONS 0 1932>
 "00000000000000000000011110001101", -- 1932 FREE #<CONS 0 1933>
 "00000000000000000000011110001110", -- 1933 FREE #<CONS 0 1934>
 "00000000000000000000011110001111", -- 1934 FREE #<CONS 0 1935>
 "00000000000000000000011110010000", -- 1935 FREE #<CONS 0 1936>
 "00000000000000000000011110010001", -- 1936 FREE #<CONS 0 1937>
 "00000000000000000000011110010010", -- 1937 FREE #<CONS 0 1938>
 "00000000000000000000011110010011", -- 1938 FREE #<CONS 0 1939>
 "00000000000000000000011110010100", -- 1939 FREE #<CONS 0 1940>
 "00000000000000000000011110010101", -- 1940 FREE #<CONS 0 1941>
 "00000000000000000000011110010110", -- 1941 FREE #<CONS 0 1942>
 "00000000000000000000011110010111", -- 1942 FREE #<CONS 0 1943>
 "00000000000000000000011110011000", -- 1943 FREE #<CONS 0 1944>
 "00000000000000000000011110011001", -- 1944 FREE #<CONS 0 1945>
 "00000000000000000000011110011010", -- 1945 FREE #<CONS 0 1946>
 "00000000000000000000011110011011", -- 1946 FREE #<CONS 0 1947>
 "00000000000000000000011110011100", -- 1947 FREE #<CONS 0 1948>
 "00000000000000000000011110011101", -- 1948 FREE #<CONS 0 1949>
 "00000000000000000000011110011110", -- 1949 FREE #<CONS 0 1950>
 "00000000000000000000011110011111", -- 1950 FREE #<CONS 0 1951>
 "00000000000000000000011110100000", -- 1951 FREE #<CONS 0 1952>
 "00000000000000000000011110100001", -- 1952 FREE #<CONS 0 1953>
 "00000000000000000000011110100010", -- 1953 FREE #<CONS 0 1954>
 "00000000000000000000011110100011", -- 1954 FREE #<CONS 0 1955>
 "00000000000000000000011110100100", -- 1955 FREE #<CONS 0 1956>
 "00000000000000000000011110100101", -- 1956 FREE #<CONS 0 1957>
 "00000000000000000000011110100110", -- 1957 FREE #<CONS 0 1958>
 "00000000000000000000011110100111", -- 1958 FREE #<CONS 0 1959>
 "00000000000000000000011110101000", -- 1959 FREE #<CONS 0 1960>
 "00000000000000000000011110101001", -- 1960 FREE #<CONS 0 1961>
 "00000000000000000000011110101010", -- 1961 FREE #<CONS 0 1962>
 "00000000000000000000011110101011", -- 1962 FREE #<CONS 0 1963>
 "00000000000000000000011110101100", -- 1963 FREE #<CONS 0 1964>
 "00000000000000000000011110101101", -- 1964 FREE #<CONS 0 1965>
 "00000000000000000000011110101110", -- 1965 FREE #<CONS 0 1966>
 "00000000000000000000011110101111", -- 1966 FREE #<CONS 0 1967>
 "00000000000000000000011110110000", -- 1967 FREE #<CONS 0 1968>
 "00000000000000000000011110110001", -- 1968 FREE #<CONS 0 1969>
 "00000000000000000000011110110010", -- 1969 FREE #<CONS 0 1970>
 "00000000000000000000011110110011", -- 1970 FREE #<CONS 0 1971>
 "00000000000000000000011110110100", -- 1971 FREE #<CONS 0 1972>
 "00000000000000000000011110110101", -- 1972 FREE #<CONS 0 1973>
 "00000000000000000000011110110110", -- 1973 FREE #<CONS 0 1974>
 "00000000000000000000011110110111", -- 1974 FREE #<CONS 0 1975>
 "00000000000000000000011110111000", -- 1975 FREE #<CONS 0 1976>
 "00000000000000000000011110111001", -- 1976 FREE #<CONS 0 1977>
 "00000000000000000000011110111010", -- 1977 FREE #<CONS 0 1978>
 "00000000000000000000011110111011", -- 1978 FREE #<CONS 0 1979>
 "00000000000000000000011110111100", -- 1979 FREE #<CONS 0 1980>
 "00000000000000000000011110111101", -- 1980 FREE #<CONS 0 1981>
 "00000000000000000000011110111110", -- 1981 FREE #<CONS 0 1982>
 "00000000000000000000011110111111", -- 1982 FREE #<CONS 0 1983>
 "00000000000000000000011111000000", -- 1983 FREE #<CONS 0 1984>
 "00000000000000000000011111000001", -- 1984 FREE #<CONS 0 1985>
 "00000000000000000000011111000010", -- 1985 FREE #<CONS 0 1986>
 "00000000000000000000011111000011", -- 1986 FREE #<CONS 0 1987>
 "00000000000000000000011111000100", -- 1987 FREE #<CONS 0 1988>
 "00000000000000000000011111000101", -- 1988 FREE #<CONS 0 1989>
 "00000000000000000000011111000110", -- 1989 FREE #<CONS 0 1990>
 "00000000000000000000011111000111", -- 1990 FREE #<CONS 0 1991>
 "00000000000000000000011111001000", -- 1991 FREE #<CONS 0 1992>
 "00000000000000000000011111001001", -- 1992 FREE #<CONS 0 1993>
 "00000000000000000000011111001010", -- 1993 FREE #<CONS 0 1994>
 "00000000000000000000011111001011", -- 1994 FREE #<CONS 0 1995>
 "00000000000000000000011111001100", -- 1995 FREE #<CONS 0 1996>
 "00000000000000000000011111001101", -- 1996 FREE #<CONS 0 1997>
 "00000000000000000000011111001110", -- 1997 FREE #<CONS 0 1998>
 "00000000000000000000011111001111", -- 1998 FREE #<CONS 0 1999>
 "00000000000000000000011111010000", -- 1999 FREE #<CONS 0 2000>
 "00000000000000000000011111010001", -- 2000 FREE #<CONS 0 2001>
 "00000000000000000000011111010010", -- 2001 FREE #<CONS 0 2002>
 "00000000000000000000011111010011", -- 2002 FREE #<CONS 0 2003>
 "00000000000000000000011111010100", -- 2003 FREE #<CONS 0 2004>
 "00000000000000000000011111010101", -- 2004 FREE #<CONS 0 2005>
 "00000000000000000000011111010110", -- 2005 FREE #<CONS 0 2006>
 "00000000000000000000011111010111", -- 2006 FREE #<CONS 0 2007>
 "00000000000000000000011111011000", -- 2007 FREE #<CONS 0 2008>
 "00000000000000000000011111011001", -- 2008 FREE #<CONS 0 2009>
 "00000000000000000000011111011010", -- 2009 FREE #<CONS 0 2010>
 "00000000000000000000011111011011", -- 2010 FREE #<CONS 0 2011>
 "00000000000000000000011111011100", -- 2011 FREE #<CONS 0 2012>
 "00000000000000000000011111011101", -- 2012 FREE #<CONS 0 2013>
 "00000000000000000000011111011110", -- 2013 FREE #<CONS 0 2014>
 "00000000000000000000011111011111", -- 2014 FREE #<CONS 0 2015>
 "00000000000000000000011111100000", -- 2015 FREE #<CONS 0 2016>
 "00000000000000000000011111100001", -- 2016 FREE #<CONS 0 2017>
 "00000000000000000000011111100010", -- 2017 FREE #<CONS 0 2018>
 "00000000000000000000011111100011", -- 2018 FREE #<CONS 0 2019>
 "00000000000000000000011111100100", -- 2019 FREE #<CONS 0 2020>
 "00000000000000000000011111100101", -- 2020 FREE #<CONS 0 2021>
 "00000000000000000000011111100110", -- 2021 FREE #<CONS 0 2022>
 "00000000000000000000011111100111", -- 2022 FREE #<CONS 0 2023>
 "00000000000000000000011111101000", -- 2023 FREE #<CONS 0 2024>
 "00000000000000000000011111101001", -- 2024 FREE #<CONS 0 2025>
 "00000000000000000000011111101010", -- 2025 FREE #<CONS 0 2026>
 "00000000000000000000011111101011", -- 2026 FREE #<CONS 0 2027>
 "00000000000000000000011111101100", -- 2027 FREE #<CONS 0 2028>
 "00000000000000000000011111101101", -- 2028 FREE #<CONS 0 2029>
 "00000000000000000000011111101110", -- 2029 FREE #<CONS 0 2030>
 "00000000000000000000011111101111", -- 2030 FREE #<CONS 0 2031>
 "00000000000000000000011111110000", -- 2031 FREE #<CONS 0 2032>
 "00000000000000000000011111110001", -- 2032 FREE #<CONS 0 2033>
 "00000000000000000000011111110010", -- 2033 FREE #<CONS 0 2034>
 "00000000000000000000011111110011", -- 2034 FREE #<CONS 0 2035>
 "00000000000000000000011111110100", -- 2035 FREE #<CONS 0 2036>
 "00000000000000000000011111110101", -- 2036 FREE #<CONS 0 2037>
 "00000000000000000000011111110110", -- 2037 FREE #<CONS 0 2038>
 "00000000000000000000011111110111", -- 2038 FREE #<CONS 0 2039>
 "00000000000000000000011111111000", -- 2039 FREE #<CONS 0 2040>
 "00000000000000000000011111111001", -- 2040 FREE #<CONS 0 2041>
 "00000000000000000000011111111010", -- 2041 FREE #<CONS 0 2042>
 "00000000000000000000011111111011", -- 2042 FREE #<CONS 0 2043>
 "00000000000000000000011111111100", -- 2043 FREE #<CONS 0 2044>
 "00000000000000000000011111111101", -- 2044 FREE #<CONS 0 2045>
 "00000000000000000000011111111110", -- 2045 FREE #<CONS 0 2046>
 "00000000000000000000011111111111", -- 2046 FREE #<CONS 0 2047>
 "00000000000000000000100000000000", -- 2047 FREE #<CONS 0 2048>
 "00000000000000000000100000000001", -- 2048 FREE #<CONS 0 2049>
 "00000000000000000000100000000010", -- 2049 FREE #<CONS 0 2050>
 "00000000000000000000100000000011", -- 2050 FREE #<CONS 0 2051>
 "00000000000000000000100000000100", -- 2051 FREE #<CONS 0 2052>
 "00000000000000000000100000000101", -- 2052 FREE #<CONS 0 2053>
 "00000000000000000000100000000110", -- 2053 FREE #<CONS 0 2054>
 "00000000000000000000100000000111", -- 2054 FREE #<CONS 0 2055>
 "00000000000000000000100000001000", -- 2055 FREE #<CONS 0 2056>
 "00000000000000000000100000001001", -- 2056 FREE #<CONS 0 2057>
 "00000000000000000000100000001010", -- 2057 FREE #<CONS 0 2058>
 "00000000000000000000100000001011", -- 2058 FREE #<CONS 0 2059>
 "00000000000000000000100000001100", -- 2059 FREE #<CONS 0 2060>
 "00000000000000000000100000001101", -- 2060 FREE #<CONS 0 2061>
 "00000000000000000000100000001110", -- 2061 FREE #<CONS 0 2062>
 "00000000000000000000100000001111", -- 2062 FREE #<CONS 0 2063>
 "00000000000000000000100000010000", -- 2063 FREE #<CONS 0 2064>
 "00000000000000000000100000010001", -- 2064 FREE #<CONS 0 2065>
 "00000000000000000000100000010010", -- 2065 FREE #<CONS 0 2066>
 "00000000000000000000100000010011", -- 2066 FREE #<CONS 0 2067>
 "00000000000000000000100000010100", -- 2067 FREE #<CONS 0 2068>
 "00000000000000000000100000010101", -- 2068 FREE #<CONS 0 2069>
 "00000000000000000000100000010110", -- 2069 FREE #<CONS 0 2070>
 "00000000000000000000100000010111", -- 2070 FREE #<CONS 0 2071>
 "00000000000000000000100000011000", -- 2071 FREE #<CONS 0 2072>
 "00000000000000000000100000011001", -- 2072 FREE #<CONS 0 2073>
 "00000000000000000000100000011010", -- 2073 FREE #<CONS 0 2074>
 "00000000000000000000100000011011", -- 2074 FREE #<CONS 0 2075>
 "00000000000000000000100000011100", -- 2075 FREE #<CONS 0 2076>
 "00000000000000000000100000011101", -- 2076 FREE #<CONS 0 2077>
 "00000000000000000000100000011110", -- 2077 FREE #<CONS 0 2078>
 "00000000000000000000100000011111", -- 2078 FREE #<CONS 0 2079>
 "00000000000000000000100000100000", -- 2079 FREE #<CONS 0 2080>
 "00000000000000000000100000100001", -- 2080 FREE #<CONS 0 2081>
 "00000000000000000000100000100010", -- 2081 FREE #<CONS 0 2082>
 "00000000000000000000100000100011", -- 2082 FREE #<CONS 0 2083>
 "00000000000000000000100000100100", -- 2083 FREE #<CONS 0 2084>
 "00000000000000000000100000100101", -- 2084 FREE #<CONS 0 2085>
 "00000000000000000000100000100110", -- 2085 FREE #<CONS 0 2086>
 "00000000000000000000100000100111", -- 2086 FREE #<CONS 0 2087>
 "00000000000000000000100000101000", -- 2087 FREE #<CONS 0 2088>
 "00000000000000000000100000101001", -- 2088 FREE #<CONS 0 2089>
 "00000000000000000000100000101010", -- 2089 FREE #<CONS 0 2090>
 "00000000000000000000100000101011", -- 2090 FREE #<CONS 0 2091>
 "00000000000000000000100000101100", -- 2091 FREE #<CONS 0 2092>
 "00000000000000000000100000101101", -- 2092 FREE #<CONS 0 2093>
 "00000000000000000000100000101110", -- 2093 FREE #<CONS 0 2094>
 "00000000000000000000100000101111", -- 2094 FREE #<CONS 0 2095>
 "00000000000000000000100000110000", -- 2095 FREE #<CONS 0 2096>
 "00000000000000000000100000110001", -- 2096 FREE #<CONS 0 2097>
 "00000000000000000000100000110010", -- 2097 FREE #<CONS 0 2098>
 "00000000000000000000100000110011", -- 2098 FREE #<CONS 0 2099>
 "00000000000000000000100000110100", -- 2099 FREE #<CONS 0 2100>
 "00000000000000000000100000110101", -- 2100 FREE #<CONS 0 2101>
 "00000000000000000000100000110110", -- 2101 FREE #<CONS 0 2102>
 "00000000000000000000100000110111", -- 2102 FREE #<CONS 0 2103>
 "00000000000000000000100000111000", -- 2103 FREE #<CONS 0 2104>
 "00000000000000000000100000111001", -- 2104 FREE #<CONS 0 2105>
 "00000000000000000000100000111010", -- 2105 FREE #<CONS 0 2106>
 "00000000000000000000100000111011", -- 2106 FREE #<CONS 0 2107>
 "00000000000000000000100000111100", -- 2107 FREE #<CONS 0 2108>
 "00000000000000000000100000111101", -- 2108 FREE #<CONS 0 2109>
 "00000000000000000000100000111110", -- 2109 FREE #<CONS 0 2110>
 "00000000000000000000100000111111", -- 2110 FREE #<CONS 0 2111>
 "00000000000000000000100001000000", -- 2111 FREE #<CONS 0 2112>
 "00000000000000000000100001000001", -- 2112 FREE #<CONS 0 2113>
 "00000000000000000000100001000010", -- 2113 FREE #<CONS 0 2114>
 "00000000000000000000100001000011", -- 2114 FREE #<CONS 0 2115>
 "00000000000000000000100001000100", -- 2115 FREE #<CONS 0 2116>
 "00000000000000000000100001000101", -- 2116 FREE #<CONS 0 2117>
 "00000000000000000000100001000110", -- 2117 FREE #<CONS 0 2118>
 "00000000000000000000100001000111", -- 2118 FREE #<CONS 0 2119>
 "00000000000000000000100001001000", -- 2119 FREE #<CONS 0 2120>
 "00000000000000000000100001001001", -- 2120 FREE #<CONS 0 2121>
 "00000000000000000000100001001010", -- 2121 FREE #<CONS 0 2122>
 "00000000000000000000100001001011", -- 2122 FREE #<CONS 0 2123>
 "00000000000000000000100001001100", -- 2123 FREE #<CONS 0 2124>
 "00000000000000000000100001001101", -- 2124 FREE #<CONS 0 2125>
 "00000000000000000000100001001110", -- 2125 FREE #<CONS 0 2126>
 "00000000000000000000100001001111", -- 2126 FREE #<CONS 0 2127>
 "00000000000000000000100001010000", -- 2127 FREE #<CONS 0 2128>
 "00000000000000000000100001010001", -- 2128 FREE #<CONS 0 2129>
 "00000000000000000000100001010010", -- 2129 FREE #<CONS 0 2130>
 "00000000000000000000100001010011", -- 2130 FREE #<CONS 0 2131>
 "00000000000000000000100001010100", -- 2131 FREE #<CONS 0 2132>
 "00000000000000000000100001010101", -- 2132 FREE #<CONS 0 2133>
 "00000000000000000000100001010110", -- 2133 FREE #<CONS 0 2134>
 "00000000000000000000100001010111", -- 2134 FREE #<CONS 0 2135>
 "00000000000000000000100001011000", -- 2135 FREE #<CONS 0 2136>
 "00000000000000000000100001011001", -- 2136 FREE #<CONS 0 2137>
 "00000000000000000000100001011010", -- 2137 FREE #<CONS 0 2138>
 "00000000000000000000100001011011", -- 2138 FREE #<CONS 0 2139>
 "00000000000000000000100001011100", -- 2139 FREE #<CONS 0 2140>
 "00000000000000000000100001011101", -- 2140 FREE #<CONS 0 2141>
 "00000000000000000000100001011110", -- 2141 FREE #<CONS 0 2142>
 "00000000000000000000100001011111", -- 2142 FREE #<CONS 0 2143>
 "00000000000000000000100001100000", -- 2143 FREE #<CONS 0 2144>
 "00000000000000000000100001100001", -- 2144 FREE #<CONS 0 2145>
 "00000000000000000000100001100010", -- 2145 FREE #<CONS 0 2146>
 "00000000000000000000100001100011", -- 2146 FREE #<CONS 0 2147>
 "00000000000000000000100001100100", -- 2147 FREE #<CONS 0 2148>
 "00000000000000000000100001100101", -- 2148 FREE #<CONS 0 2149>
 "00000000000000000000100001100110", -- 2149 FREE #<CONS 0 2150>
 "00000000000000000000100001100111", -- 2150 FREE #<CONS 0 2151>
 "00000000000000000000100001101000", -- 2151 FREE #<CONS 0 2152>
 "00000000000000000000100001101001", -- 2152 FREE #<CONS 0 2153>
 "00000000000000000000100001101010", -- 2153 FREE #<CONS 0 2154>
 "00000000000000000000100001101011", -- 2154 FREE #<CONS 0 2155>
 "00000000000000000000100001101100", -- 2155 FREE #<CONS 0 2156>
 "00000000000000000000100001101101", -- 2156 FREE #<CONS 0 2157>
 "00000000000000000000100001101110", -- 2157 FREE #<CONS 0 2158>
 "00000000000000000000100001101111", -- 2158 FREE #<CONS 0 2159>
 "00000000000000000000100001110000", -- 2159 FREE #<CONS 0 2160>
 "00000000000000000000100001110001", -- 2160 FREE #<CONS 0 2161>
 "00000000000000000000100001110010", -- 2161 FREE #<CONS 0 2162>
 "00000000000000000000100001110011", -- 2162 FREE #<CONS 0 2163>
 "00000000000000000000100001110100", -- 2163 FREE #<CONS 0 2164>
 "00000000000000000000100001110101", -- 2164 FREE #<CONS 0 2165>
 "00000000000000000000100001110110", -- 2165 FREE #<CONS 0 2166>
 "00000000000000000000100001110111", -- 2166 FREE #<CONS 0 2167>
 "00000000000000000000100001111000", -- 2167 FREE #<CONS 0 2168>
 "00000000000000000000100001111001", -- 2168 FREE #<CONS 0 2169>
 "00000000000000000000100001111010", -- 2169 FREE #<CONS 0 2170>
 "00000000000000000000100001111011", -- 2170 FREE #<CONS 0 2171>
 "00000000000000000000100001111100", -- 2171 FREE #<CONS 0 2172>
 "00000000000000000000100001111101", -- 2172 FREE #<CONS 0 2173>
 "00000000000000000000100001111110", -- 2173 FREE #<CONS 0 2174>
 "00000000000000000000100001111111", -- 2174 FREE #<CONS 0 2175>
 "00000000000000000000100010000000", -- 2175 FREE #<CONS 0 2176>
 "00000000000000000000100010000001", -- 2176 FREE #<CONS 0 2177>
 "00000000000000000000100010000010", -- 2177 FREE #<CONS 0 2178>
 "00000000000000000000100010000011", -- 2178 FREE #<CONS 0 2179>
 "00000000000000000000100010000100", -- 2179 FREE #<CONS 0 2180>
 "00000000000000000000100010000101", -- 2180 FREE #<CONS 0 2181>
 "00000000000000000000100010000110", -- 2181 FREE #<CONS 0 2182>
 "00000000000000000000100010000111", -- 2182 FREE #<CONS 0 2183>
 "00000000000000000000100010001000", -- 2183 FREE #<CONS 0 2184>
 "00000000000000000000100010001001", -- 2184 FREE #<CONS 0 2185>
 "00000000000000000000100010001010", -- 2185 FREE #<CONS 0 2186>
 "00000000000000000000100010001011", -- 2186 FREE #<CONS 0 2187>
 "00000000000000000000100010001100", -- 2187 FREE #<CONS 0 2188>
 "00000000000000000000100010001101", -- 2188 FREE #<CONS 0 2189>
 "00000000000000000000100010001110", -- 2189 FREE #<CONS 0 2190>
 "00000000000000000000100010001111", -- 2190 FREE #<CONS 0 2191>
 "00000000000000000000100010010000", -- 2191 FREE #<CONS 0 2192>
 "00000000000000000000100010010001", -- 2192 FREE #<CONS 0 2193>
 "00000000000000000000100010010010", -- 2193 FREE #<CONS 0 2194>
 "00000000000000000000100010010011", -- 2194 FREE #<CONS 0 2195>
 "00000000000000000000100010010100", -- 2195 FREE #<CONS 0 2196>
 "00000000000000000000100010010101", -- 2196 FREE #<CONS 0 2197>
 "00000000000000000000100010010110", -- 2197 FREE #<CONS 0 2198>
 "00000000000000000000100010010111", -- 2198 FREE #<CONS 0 2199>
 "00000000000000000000100010011000", -- 2199 FREE #<CONS 0 2200>
 "00000000000000000000100010011001", -- 2200 FREE #<CONS 0 2201>
 "00000000000000000000100010011010", -- 2201 FREE #<CONS 0 2202>
 "00000000000000000000100010011011", -- 2202 FREE #<CONS 0 2203>
 "00000000000000000000100010011100", -- 2203 FREE #<CONS 0 2204>
 "00000000000000000000100010011101", -- 2204 FREE #<CONS 0 2205>
 "00000000000000000000100010011110", -- 2205 FREE #<CONS 0 2206>
 "00000000000000000000100010011111", -- 2206 FREE #<CONS 0 2207>
 "00000000000000000000100010100000", -- 2207 FREE #<CONS 0 2208>
 "00000000000000000000100010100001", -- 2208 FREE #<CONS 0 2209>
 "00000000000000000000100010100010", -- 2209 FREE #<CONS 0 2210>
 "00000000000000000000100010100011", -- 2210 FREE #<CONS 0 2211>
 "00000000000000000000100010100100", -- 2211 FREE #<CONS 0 2212>
 "00000000000000000000100010100101", -- 2212 FREE #<CONS 0 2213>
 "00000000000000000000100010100110", -- 2213 FREE #<CONS 0 2214>
 "00000000000000000000100010100111", -- 2214 FREE #<CONS 0 2215>
 "00000000000000000000100010101000", -- 2215 FREE #<CONS 0 2216>
 "00000000000000000000100010101001", -- 2216 FREE #<CONS 0 2217>
 "00000000000000000000100010101010", -- 2217 FREE #<CONS 0 2218>
 "00000000000000000000100010101011", -- 2218 FREE #<CONS 0 2219>
 "00000000000000000000100010101100", -- 2219 FREE #<CONS 0 2220>
 "00000000000000000000100010101101", -- 2220 FREE #<CONS 0 2221>
 "00000000000000000000100010101110", -- 2221 FREE #<CONS 0 2222>
 "00000000000000000000100010101111", -- 2222 FREE #<CONS 0 2223>
 "00000000000000000000100010110000", -- 2223 FREE #<CONS 0 2224>
 "00000000000000000000100010110001", -- 2224 FREE #<CONS 0 2225>
 "00000000000000000000100010110010", -- 2225 FREE #<CONS 0 2226>
 "00000000000000000000100010110011", -- 2226 FREE #<CONS 0 2227>
 "00000000000000000000100010110100", -- 2227 FREE #<CONS 0 2228>
 "00000000000000000000100010110101", -- 2228 FREE #<CONS 0 2229>
 "00000000000000000000100010110110", -- 2229 FREE #<CONS 0 2230>
 "00000000000000000000100010110111", -- 2230 FREE #<CONS 0 2231>
 "00000000000000000000100010111000", -- 2231 FREE #<CONS 0 2232>
 "00000000000000000000100010111001", -- 2232 FREE #<CONS 0 2233>
 "00000000000000000000100010111010", -- 2233 FREE #<CONS 0 2234>
 "00000000000000000000100010111011", -- 2234 FREE #<CONS 0 2235>
 "00000000000000000000100010111100", -- 2235 FREE #<CONS 0 2236>
 "00000000000000000000100010111101", -- 2236 FREE #<CONS 0 2237>
 "00000000000000000000100010111110", -- 2237 FREE #<CONS 0 2238>
 "00000000000000000000100010111111", -- 2238 FREE #<CONS 0 2239>
 "00000000000000000000100011000000", -- 2239 FREE #<CONS 0 2240>
 "00000000000000000000100011000001", -- 2240 FREE #<CONS 0 2241>
 "00000000000000000000100011000010", -- 2241 FREE #<CONS 0 2242>
 "00000000000000000000100011000011", -- 2242 FREE #<CONS 0 2243>
 "00000000000000000000100011000100", -- 2243 FREE #<CONS 0 2244>
 "00000000000000000000100011000101", -- 2244 FREE #<CONS 0 2245>
 "00000000000000000000100011000110", -- 2245 FREE #<CONS 0 2246>
 "00000000000000000000100011000111", -- 2246 FREE #<CONS 0 2247>
 "00000000000000000000100011001000", -- 2247 FREE #<CONS 0 2248>
 "00000000000000000000100011001001", -- 2248 FREE #<CONS 0 2249>
 "00000000000000000000100011001010", -- 2249 FREE #<CONS 0 2250>
 "00000000000000000000100011001011", -- 2250 FREE #<CONS 0 2251>
 "00000000000000000000100011001100", -- 2251 FREE #<CONS 0 2252>
 "00000000000000000000100011001101", -- 2252 FREE #<CONS 0 2253>
 "00000000000000000000100011001110", -- 2253 FREE #<CONS 0 2254>
 "00000000000000000000100011001111", -- 2254 FREE #<CONS 0 2255>
 "00000000000000000000100011010000", -- 2255 FREE #<CONS 0 2256>
 "00000000000000000000100011010001", -- 2256 FREE #<CONS 0 2257>
 "00000000000000000000100011010010", -- 2257 FREE #<CONS 0 2258>
 "00000000000000000000100011010011", -- 2258 FREE #<CONS 0 2259>
 "00000000000000000000100011010100", -- 2259 FREE #<CONS 0 2260>
 "00000000000000000000100011010101", -- 2260 FREE #<CONS 0 2261>
 "00000000000000000000100011010110", -- 2261 FREE #<CONS 0 2262>
 "00000000000000000000100011010111", -- 2262 FREE #<CONS 0 2263>
 "00000000000000000000100011011000", -- 2263 FREE #<CONS 0 2264>
 "00000000000000000000100011011001", -- 2264 FREE #<CONS 0 2265>
 "00000000000000000000100011011010", -- 2265 FREE #<CONS 0 2266>
 "00000000000000000000100011011011", -- 2266 FREE #<CONS 0 2267>
 "00000000000000000000100011011100", -- 2267 FREE #<CONS 0 2268>
 "00000000000000000000100011011101", -- 2268 FREE #<CONS 0 2269>
 "00000000000000000000100011011110", -- 2269 FREE #<CONS 0 2270>
 "00000000000000000000100011011111", -- 2270 FREE #<CONS 0 2271>
 "00000000000000000000100011100000", -- 2271 FREE #<CONS 0 2272>
 "00000000000000000000100011100001", -- 2272 FREE #<CONS 0 2273>
 "00000000000000000000100011100010", -- 2273 FREE #<CONS 0 2274>
 "00000000000000000000100011100011", -- 2274 FREE #<CONS 0 2275>
 "00000000000000000000100011100100", -- 2275 FREE #<CONS 0 2276>
 "00000000000000000000100011100101", -- 2276 FREE #<CONS 0 2277>
 "00000000000000000000100011100110", -- 2277 FREE #<CONS 0 2278>
 "00000000000000000000100011100111", -- 2278 FREE #<CONS 0 2279>
 "00000000000000000000100011101000", -- 2279 FREE #<CONS 0 2280>
 "00000000000000000000100011101001", -- 2280 FREE #<CONS 0 2281>
 "00000000000000000000100011101010", -- 2281 FREE #<CONS 0 2282>
 "00000000000000000000100011101011", -- 2282 FREE #<CONS 0 2283>
 "00000000000000000000100011101100", -- 2283 FREE #<CONS 0 2284>
 "00000000000000000000100011101101", -- 2284 FREE #<CONS 0 2285>
 "00000000000000000000100011101110", -- 2285 FREE #<CONS 0 2286>
 "00000000000000000000100011101111", -- 2286 FREE #<CONS 0 2287>
 "00000000000000000000100011110000", -- 2287 FREE #<CONS 0 2288>
 "00000000000000000000100011110001", -- 2288 FREE #<CONS 0 2289>
 "00000000000000000000100011110010", -- 2289 FREE #<CONS 0 2290>
 "00000000000000000000100011110011", -- 2290 FREE #<CONS 0 2291>
 "00000000000000000000100011110100", -- 2291 FREE #<CONS 0 2292>
 "00000000000000000000100011110101", -- 2292 FREE #<CONS 0 2293>
 "00000000000000000000100011110110", -- 2293 FREE #<CONS 0 2294>
 "00000000000000000000100011110111", -- 2294 FREE #<CONS 0 2295>
 "00000000000000000000100011111000", -- 2295 FREE #<CONS 0 2296>
 "00000000000000000000100011111001", -- 2296 FREE #<CONS 0 2297>
 "00000000000000000000100011111010", -- 2297 FREE #<CONS 0 2298>
 "00000000000000000000100011111011", -- 2298 FREE #<CONS 0 2299>
 "00000000000000000000100011111100", -- 2299 FREE #<CONS 0 2300>
 "00000000000000000000100011111101", -- 2300 FREE #<CONS 0 2301>
 "00000000000000000000100011111110", -- 2301 FREE #<CONS 0 2302>
 "00000000000000000000100011111111", -- 2302 FREE #<CONS 0 2303>
 "00000000000000000000100100000000", -- 2303 FREE #<CONS 0 2304>
 "00000000000000000000100100000001", -- 2304 FREE #<CONS 0 2305>
 "00000000000000000000100100000010", -- 2305 FREE #<CONS 0 2306>
 "00000000000000000000100100000011", -- 2306 FREE #<CONS 0 2307>
 "00000000000000000000100100000100", -- 2307 FREE #<CONS 0 2308>
 "00000000000000000000100100000101", -- 2308 FREE #<CONS 0 2309>
 "00000000000000000000100100000110", -- 2309 FREE #<CONS 0 2310>
 "00000000000000000000100100000111", -- 2310 FREE #<CONS 0 2311>
 "00000000000000000000100100001000", -- 2311 FREE #<CONS 0 2312>
 "00000000000000000000100100001001", -- 2312 FREE #<CONS 0 2313>
 "00000000000000000000100100001010", -- 2313 FREE #<CONS 0 2314>
 "00000000000000000000100100001011", -- 2314 FREE #<CONS 0 2315>
 "00000000000000000000100100001100", -- 2315 FREE #<CONS 0 2316>
 "00000000000000000000100100001101", -- 2316 FREE #<CONS 0 2317>
 "00000000000000000000100100001110", -- 2317 FREE #<CONS 0 2318>
 "00000000000000000000100100001111", -- 2318 FREE #<CONS 0 2319>
 "00000000000000000000100100010000", -- 2319 FREE #<CONS 0 2320>
 "00000000000000000000100100010001", -- 2320 FREE #<CONS 0 2321>
 "00000000000000000000100100010010", -- 2321 FREE #<CONS 0 2322>
 "00000000000000000000100100010011", -- 2322 FREE #<CONS 0 2323>
 "00000000000000000000100100010100", -- 2323 FREE #<CONS 0 2324>
 "00000000000000000000100100010101", -- 2324 FREE #<CONS 0 2325>
 "00000000000000000000100100010110", -- 2325 FREE #<CONS 0 2326>
 "00000000000000000000100100010111", -- 2326 FREE #<CONS 0 2327>
 "00000000000000000000100100011000", -- 2327 FREE #<CONS 0 2328>
 "00000000000000000000100100011001", -- 2328 FREE #<CONS 0 2329>
 "00000000000000000000100100011010", -- 2329 FREE #<CONS 0 2330>
 "00000000000000000000100100011011", -- 2330 FREE #<CONS 0 2331>
 "00000000000000000000100100011100", -- 2331 FREE #<CONS 0 2332>
 "00000000000000000000100100011101", -- 2332 FREE #<CONS 0 2333>
 "00000000000000000000100100011110", -- 2333 FREE #<CONS 0 2334>
 "00000000000000000000100100011111", -- 2334 FREE #<CONS 0 2335>
 "00000000000000000000100100100000", -- 2335 FREE #<CONS 0 2336>
 "00000000000000000000100100100001", -- 2336 FREE #<CONS 0 2337>
 "00000000000000000000100100100010", -- 2337 FREE #<CONS 0 2338>
 "00000000000000000000100100100011", -- 2338 FREE #<CONS 0 2339>
 "00000000000000000000100100100100", -- 2339 FREE #<CONS 0 2340>
 "00000000000000000000100100100101", -- 2340 FREE #<CONS 0 2341>
 "00000000000000000000100100100110", -- 2341 FREE #<CONS 0 2342>
 "00000000000000000000100100100111", -- 2342 FREE #<CONS 0 2343>
 "00000000000000000000100100101000", -- 2343 FREE #<CONS 0 2344>
 "00000000000000000000100100101001", -- 2344 FREE #<CONS 0 2345>
 "00000000000000000000100100101010", -- 2345 FREE #<CONS 0 2346>
 "00000000000000000000100100101011", -- 2346 FREE #<CONS 0 2347>
 "00000000000000000000100100101100", -- 2347 FREE #<CONS 0 2348>
 "00000000000000000000100100101101", -- 2348 FREE #<CONS 0 2349>
 "00000000000000000000100100101110", -- 2349 FREE #<CONS 0 2350>
 "00000000000000000000100100101111", -- 2350 FREE #<CONS 0 2351>
 "00000000000000000000100100110000", -- 2351 FREE #<CONS 0 2352>
 "00000000000000000000100100110001", -- 2352 FREE #<CONS 0 2353>
 "00000000000000000000100100110010", -- 2353 FREE #<CONS 0 2354>
 "00000000000000000000100100110011", -- 2354 FREE #<CONS 0 2355>
 "00000000000000000000100100110100", -- 2355 FREE #<CONS 0 2356>
 "00000000000000000000100100110101", -- 2356 FREE #<CONS 0 2357>
 "00000000000000000000100100110110", -- 2357 FREE #<CONS 0 2358>
 "00000000000000000000100100110111", -- 2358 FREE #<CONS 0 2359>
 "00000000000000000000100100111000", -- 2359 FREE #<CONS 0 2360>
 "00000000000000000000100100111001", -- 2360 FREE #<CONS 0 2361>
 "00000000000000000000100100111010", -- 2361 FREE #<CONS 0 2362>
 "00000000000000000000100100111011", -- 2362 FREE #<CONS 0 2363>
 "00000000000000000000100100111100", -- 2363 FREE #<CONS 0 2364>
 "00000000000000000000100100111101", -- 2364 FREE #<CONS 0 2365>
 "00000000000000000000100100111110", -- 2365 FREE #<CONS 0 2366>
 "00000000000000000000100100111111", -- 2366 FREE #<CONS 0 2367>
 "00000000000000000000100101000000", -- 2367 FREE #<CONS 0 2368>
 "00000000000000000000100101000001", -- 2368 FREE #<CONS 0 2369>
 "00000000000000000000100101000010", -- 2369 FREE #<CONS 0 2370>
 "00000000000000000000100101000011", -- 2370 FREE #<CONS 0 2371>
 "00000000000000000000100101000100", -- 2371 FREE #<CONS 0 2372>
 "00000000000000000000100101000101", -- 2372 FREE #<CONS 0 2373>
 "00000000000000000000100101000110", -- 2373 FREE #<CONS 0 2374>
 "00000000000000000000100101000111", -- 2374 FREE #<CONS 0 2375>
 "00000000000000000000100101001000", -- 2375 FREE #<CONS 0 2376>
 "00000000000000000000100101001001", -- 2376 FREE #<CONS 0 2377>
 "00000000000000000000100101001010", -- 2377 FREE #<CONS 0 2378>
 "00000000000000000000100101001011", -- 2378 FREE #<CONS 0 2379>
 "00000000000000000000100101001100", -- 2379 FREE #<CONS 0 2380>
 "00000000000000000000100101001101", -- 2380 FREE #<CONS 0 2381>
 "00000000000000000000100101001110", -- 2381 FREE #<CONS 0 2382>
 "00000000000000000000100101001111", -- 2382 FREE #<CONS 0 2383>
 "00000000000000000000100101010000", -- 2383 FREE #<CONS 0 2384>
 "00000000000000000000100101010001", -- 2384 FREE #<CONS 0 2385>
 "00000000000000000000100101010010", -- 2385 FREE #<CONS 0 2386>
 "00000000000000000000100101010011", -- 2386 FREE #<CONS 0 2387>
 "00000000000000000000100101010100", -- 2387 FREE #<CONS 0 2388>
 "00000000000000000000100101010101", -- 2388 FREE #<CONS 0 2389>
 "00000000000000000000100101010110", -- 2389 FREE #<CONS 0 2390>
 "00000000000000000000100101010111", -- 2390 FREE #<CONS 0 2391>
 "00000000000000000000100101011000", -- 2391 FREE #<CONS 0 2392>
 "00000000000000000000100101011001", -- 2392 FREE #<CONS 0 2393>
 "00000000000000000000100101011010", -- 2393 FREE #<CONS 0 2394>
 "00000000000000000000100101011011", -- 2394 FREE #<CONS 0 2395>
 "00000000000000000000100101011100", -- 2395 FREE #<CONS 0 2396>
 "00000000000000000000100101011101", -- 2396 FREE #<CONS 0 2397>
 "00000000000000000000100101011110", -- 2397 FREE #<CONS 0 2398>
 "00000000000000000000100101011111", -- 2398 FREE #<CONS 0 2399>
 "00000000000000000000100101100000", -- 2399 FREE #<CONS 0 2400>
 "00000000000000000000100101100001", -- 2400 FREE #<CONS 0 2401>
 "00000000000000000000100101100010", -- 2401 FREE #<CONS 0 2402>
 "00000000000000000000100101100011", -- 2402 FREE #<CONS 0 2403>
 "00000000000000000000100101100100", -- 2403 FREE #<CONS 0 2404>
 "00000000000000000000100101100101", -- 2404 FREE #<CONS 0 2405>
 "00000000000000000000100101100110", -- 2405 FREE #<CONS 0 2406>
 "00000000000000000000100101100111", -- 2406 FREE #<CONS 0 2407>
 "00000000000000000000100101101000", -- 2407 FREE #<CONS 0 2408>
 "00000000000000000000100101101001", -- 2408 FREE #<CONS 0 2409>
 "00000000000000000000100101101010", -- 2409 FREE #<CONS 0 2410>
 "00000000000000000000100101101011", -- 2410 FREE #<CONS 0 2411>
 "00000000000000000000100101101100", -- 2411 FREE #<CONS 0 2412>
 "00000000000000000000100101101101", -- 2412 FREE #<CONS 0 2413>
 "00000000000000000000100101101110", -- 2413 FREE #<CONS 0 2414>
 "00000000000000000000100101101111", -- 2414 FREE #<CONS 0 2415>
 "00000000000000000000100101110000", -- 2415 FREE #<CONS 0 2416>
 "00000000000000000000100101110001", -- 2416 FREE #<CONS 0 2417>
 "00000000000000000000100101110010", -- 2417 FREE #<CONS 0 2418>
 "00000000000000000000100101110011", -- 2418 FREE #<CONS 0 2419>
 "00000000000000000000100101110100", -- 2419 FREE #<CONS 0 2420>
 "00000000000000000000100101110101", -- 2420 FREE #<CONS 0 2421>
 "00000000000000000000100101110110", -- 2421 FREE #<CONS 0 2422>
 "00000000000000000000100101110111", -- 2422 FREE #<CONS 0 2423>
 "00000000000000000000100101111000", -- 2423 FREE #<CONS 0 2424>
 "00000000000000000000100101111001", -- 2424 FREE #<CONS 0 2425>
 "00000000000000000000100101111010", -- 2425 FREE #<CONS 0 2426>
 "00000000000000000000100101111011", -- 2426 FREE #<CONS 0 2427>
 "00000000000000000000100101111100", -- 2427 FREE #<CONS 0 2428>
 "00000000000000000000100101111101", -- 2428 FREE #<CONS 0 2429>
 "00000000000000000000100101111110", -- 2429 FREE #<CONS 0 2430>
 "00000000000000000000100101111111", -- 2430 FREE #<CONS 0 2431>
 "00000000000000000000100110000000", -- 2431 FREE #<CONS 0 2432>
 "00000000000000000000100110000001", -- 2432 FREE #<CONS 0 2433>
 "00000000000000000000100110000010", -- 2433 FREE #<CONS 0 2434>
 "00000000000000000000100110000011", -- 2434 FREE #<CONS 0 2435>
 "00000000000000000000100110000100", -- 2435 FREE #<CONS 0 2436>
 "00000000000000000000100110000101", -- 2436 FREE #<CONS 0 2437>
 "00000000000000000000100110000110", -- 2437 FREE #<CONS 0 2438>
 "00000000000000000000100110000111", -- 2438 FREE #<CONS 0 2439>
 "00000000000000000000100110001000", -- 2439 FREE #<CONS 0 2440>
 "00000000000000000000100110001001", -- 2440 FREE #<CONS 0 2441>
 "00000000000000000000100110001010", -- 2441 FREE #<CONS 0 2442>
 "00000000000000000000100110001011", -- 2442 FREE #<CONS 0 2443>
 "00000000000000000000100110001100", -- 2443 FREE #<CONS 0 2444>
 "00000000000000000000100110001101", -- 2444 FREE #<CONS 0 2445>
 "00000000000000000000100110001110", -- 2445 FREE #<CONS 0 2446>
 "00000000000000000000100110001111", -- 2446 FREE #<CONS 0 2447>
 "00000000000000000000100110010000", -- 2447 FREE #<CONS 0 2448>
 "00000000000000000000100110010001", -- 2448 FREE #<CONS 0 2449>
 "00000000000000000000100110010010", -- 2449 FREE #<CONS 0 2450>
 "00000000000000000000100110010011", -- 2450 FREE #<CONS 0 2451>
 "00000000000000000000100110010100", -- 2451 FREE #<CONS 0 2452>
 "00000000000000000000100110010101", -- 2452 FREE #<CONS 0 2453>
 "00000000000000000000100110010110", -- 2453 FREE #<CONS 0 2454>
 "00000000000000000000100110010111", -- 2454 FREE #<CONS 0 2455>
 "00000000000000000000100110011000", -- 2455 FREE #<CONS 0 2456>
 "00000000000000000000100110011001", -- 2456 FREE #<CONS 0 2457>
 "00000000000000000000100110011010", -- 2457 FREE #<CONS 0 2458>
 "00000000000000000000100110011011", -- 2458 FREE #<CONS 0 2459>
 "00000000000000000000100110011100", -- 2459 FREE #<CONS 0 2460>
 "00000000000000000000100110011101", -- 2460 FREE #<CONS 0 2461>
 "00000000000000000000100110011110", -- 2461 FREE #<CONS 0 2462>
 "00000000000000000000100110011111", -- 2462 FREE #<CONS 0 2463>
 "00000000000000000000100110100000", -- 2463 FREE #<CONS 0 2464>
 "00000000000000000000100110100001", -- 2464 FREE #<CONS 0 2465>
 "00000000000000000000100110100010", -- 2465 FREE #<CONS 0 2466>
 "00000000000000000000100110100011", -- 2466 FREE #<CONS 0 2467>
 "00000000000000000000100110100100", -- 2467 FREE #<CONS 0 2468>
 "00000000000000000000100110100101", -- 2468 FREE #<CONS 0 2469>
 "00000000000000000000100110100110", -- 2469 FREE #<CONS 0 2470>
 "00000000000000000000100110100111", -- 2470 FREE #<CONS 0 2471>
 "00000000000000000000100110101000", -- 2471 FREE #<CONS 0 2472>
 "00000000000000000000100110101001", -- 2472 FREE #<CONS 0 2473>
 "00000000000000000000100110101010", -- 2473 FREE #<CONS 0 2474>
 "00000000000000000000100110101011", -- 2474 FREE #<CONS 0 2475>
 "00000000000000000000100110101100", -- 2475 FREE #<CONS 0 2476>
 "00000000000000000000100110101101", -- 2476 FREE #<CONS 0 2477>
 "00000000000000000000100110101110", -- 2477 FREE #<CONS 0 2478>
 "00000000000000000000100110101111", -- 2478 FREE #<CONS 0 2479>
 "00000000000000000000100110110000", -- 2479 FREE #<CONS 0 2480>
 "00000000000000000000100110110001", -- 2480 FREE #<CONS 0 2481>
 "00000000000000000000100110110010", -- 2481 FREE #<CONS 0 2482>
 "00000000000000000000100110110011", -- 2482 FREE #<CONS 0 2483>
 "00000000000000000000100110110100", -- 2483 FREE #<CONS 0 2484>
 "00000000000000000000100110110101", -- 2484 FREE #<CONS 0 2485>
 "00000000000000000000100110110110", -- 2485 FREE #<CONS 0 2486>
 "00000000000000000000100110110111", -- 2486 FREE #<CONS 0 2487>
 "00000000000000000000100110111000", -- 2487 FREE #<CONS 0 2488>
 "00000000000000000000100110111001", -- 2488 FREE #<CONS 0 2489>
 "00000000000000000000100110111010", -- 2489 FREE #<CONS 0 2490>
 "00000000000000000000100110111011", -- 2490 FREE #<CONS 0 2491>
 "00000000000000000000100110111100", -- 2491 FREE #<CONS 0 2492>
 "00000000000000000000100110111101", -- 2492 FREE #<CONS 0 2493>
 "00000000000000000000100110111110", -- 2493 FREE #<CONS 0 2494>
 "00000000000000000000100110111111", -- 2494 FREE #<CONS 0 2495>
 "00000000000000000000100111000000", -- 2495 FREE #<CONS 0 2496>
 "00000000000000000000100111000001", -- 2496 FREE #<CONS 0 2497>
 "00000000000000000000100111000010", -- 2497 FREE #<CONS 0 2498>
 "00000000000000000000100111000011", -- 2498 FREE #<CONS 0 2499>
 "00000000000000000000100111000100", -- 2499 FREE #<CONS 0 2500>
 "00000000000000000000100111000101", -- 2500 FREE #<CONS 0 2501>
 "00000000000000000000100111000110", -- 2501 FREE #<CONS 0 2502>
 "00000000000000000000100111000111", -- 2502 FREE #<CONS 0 2503>
 "00000000000000000000100111001000", -- 2503 FREE #<CONS 0 2504>
 "00000000000000000000100111001001", -- 2504 FREE #<CONS 0 2505>
 "00000000000000000000100111001010", -- 2505 FREE #<CONS 0 2506>
 "00000000000000000000100111001011", -- 2506 FREE #<CONS 0 2507>
 "00000000000000000000100111001100", -- 2507 FREE #<CONS 0 2508>
 "00000000000000000000100111001101", -- 2508 FREE #<CONS 0 2509>
 "00000000000000000000100111001110", -- 2509 FREE #<CONS 0 2510>
 "00000000000000000000100111001111", -- 2510 FREE #<CONS 0 2511>
 "00000000000000000000100111010000", -- 2511 FREE #<CONS 0 2512>
 "00000000000000000000100111010001", -- 2512 FREE #<CONS 0 2513>
 "00000000000000000000100111010010", -- 2513 FREE #<CONS 0 2514>
 "00000000000000000000100111010011", -- 2514 FREE #<CONS 0 2515>
 "00000000000000000000100111010100", -- 2515 FREE #<CONS 0 2516>
 "00000000000000000000100111010101", -- 2516 FREE #<CONS 0 2517>
 "00000000000000000000100111010110", -- 2517 FREE #<CONS 0 2518>
 "00000000000000000000100111010111", -- 2518 FREE #<CONS 0 2519>
 "00000000000000000000100111011000", -- 2519 FREE #<CONS 0 2520>
 "00000000000000000000100111011001", -- 2520 FREE #<CONS 0 2521>
 "00000000000000000000100111011010", -- 2521 FREE #<CONS 0 2522>
 "00000000000000000000100111011011", -- 2522 FREE #<CONS 0 2523>
 "00000000000000000000100111011100", -- 2523 FREE #<CONS 0 2524>
 "00000000000000000000100111011101", -- 2524 FREE #<CONS 0 2525>
 "00000000000000000000100111011110", -- 2525 FREE #<CONS 0 2526>
 "00000000000000000000100111011111", -- 2526 FREE #<CONS 0 2527>
 "00000000000000000000100111100000", -- 2527 FREE #<CONS 0 2528>
 "00000000000000000000100111100001", -- 2528 FREE #<CONS 0 2529>
 "00000000000000000000100111100010", -- 2529 FREE #<CONS 0 2530>
 "00000000000000000000100111100011", -- 2530 FREE #<CONS 0 2531>
 "00000000000000000000100111100100", -- 2531 FREE #<CONS 0 2532>
 "00000000000000000000100111100101", -- 2532 FREE #<CONS 0 2533>
 "00000000000000000000100111100110", -- 2533 FREE #<CONS 0 2534>
 "00000000000000000000100111100111", -- 2534 FREE #<CONS 0 2535>
 "00000000000000000000100111101000", -- 2535 FREE #<CONS 0 2536>
 "00000000000000000000100111101001", -- 2536 FREE #<CONS 0 2537>
 "00000000000000000000100111101010", -- 2537 FREE #<CONS 0 2538>
 "00000000000000000000100111101011", -- 2538 FREE #<CONS 0 2539>
 "00000000000000000000100111101100", -- 2539 FREE #<CONS 0 2540>
 "00000000000000000000100111101101", -- 2540 FREE #<CONS 0 2541>
 "00000000000000000000100111101110", -- 2541 FREE #<CONS 0 2542>
 "00000000000000000000100111101111", -- 2542 FREE #<CONS 0 2543>
 "00000000000000000000100111110000", -- 2543 FREE #<CONS 0 2544>
 "00000000000000000000100111110001", -- 2544 FREE #<CONS 0 2545>
 "00000000000000000000100111110010", -- 2545 FREE #<CONS 0 2546>
 "00000000000000000000100111110011", -- 2546 FREE #<CONS 0 2547>
 "00000000000000000000100111110100", -- 2547 FREE #<CONS 0 2548>
 "00000000000000000000100111110101", -- 2548 FREE #<CONS 0 2549>
 "00000000000000000000100111110110", -- 2549 FREE #<CONS 0 2550>
 "00000000000000000000100111110111", -- 2550 FREE #<CONS 0 2551>
 "00000000000000000000100111111000", -- 2551 FREE #<CONS 0 2552>
 "00000000000000000000100111111001", -- 2552 FREE #<CONS 0 2553>
 "00000000000000000000100111111010", -- 2553 FREE #<CONS 0 2554>
 "00000000000000000000100111111011", -- 2554 FREE #<CONS 0 2555>
 "00000000000000000000100111111100", -- 2555 FREE #<CONS 0 2556>
 "00000000000000000000100111111101", -- 2556 FREE #<CONS 0 2557>
 "00000000000000000000100111111110", -- 2557 FREE #<CONS 0 2558>
 "00000000000000000000100111111111", -- 2558 FREE #<CONS 0 2559>
 "00000000000000000000101000000000", -- 2559 FREE #<CONS 0 2560>
 "00000000000000000000101000000001", -- 2560 FREE #<CONS 0 2561>
 "00000000000000000000101000000010", -- 2561 FREE #<CONS 0 2562>
 "00000000000000000000101000000011", -- 2562 FREE #<CONS 0 2563>
 "00000000000000000000101000000100", -- 2563 FREE #<CONS 0 2564>
 "00000000000000000000101000000101", -- 2564 FREE #<CONS 0 2565>
 "00000000000000000000101000000110", -- 2565 FREE #<CONS 0 2566>
 "00000000000000000000101000000111", -- 2566 FREE #<CONS 0 2567>
 "00000000000000000000101000001000", -- 2567 FREE #<CONS 0 2568>
 "00000000000000000000101000001001", -- 2568 FREE #<CONS 0 2569>
 "00000000000000000000101000001010", -- 2569 FREE #<CONS 0 2570>
 "00000000000000000000101000001011", -- 2570 FREE #<CONS 0 2571>
 "00000000000000000000101000001100", -- 2571 FREE #<CONS 0 2572>
 "00000000000000000000101000001101", -- 2572 FREE #<CONS 0 2573>
 "00000000000000000000101000001110", -- 2573 FREE #<CONS 0 2574>
 "00000000000000000000101000001111", -- 2574 FREE #<CONS 0 2575>
 "00000000000000000000101000010000", -- 2575 FREE #<CONS 0 2576>
 "00000000000000000000101000010001", -- 2576 FREE #<CONS 0 2577>
 "00000000000000000000101000010010", -- 2577 FREE #<CONS 0 2578>
 "00000000000000000000101000010011", -- 2578 FREE #<CONS 0 2579>
 "00000000000000000000101000010100", -- 2579 FREE #<CONS 0 2580>
 "00000000000000000000101000010101", -- 2580 FREE #<CONS 0 2581>
 "00000000000000000000101000010110", -- 2581 FREE #<CONS 0 2582>
 "00000000000000000000101000010111", -- 2582 FREE #<CONS 0 2583>
 "00000000000000000000101000011000", -- 2583 FREE #<CONS 0 2584>
 "00000000000000000000101000011001", -- 2584 FREE #<CONS 0 2585>
 "00000000000000000000101000011010", -- 2585 FREE #<CONS 0 2586>
 "00000000000000000000101000011011", -- 2586 FREE #<CONS 0 2587>
 "00000000000000000000101000011100", -- 2587 FREE #<CONS 0 2588>
 "00000000000000000000101000011101", -- 2588 FREE #<CONS 0 2589>
 "00000000000000000000101000011110", -- 2589 FREE #<CONS 0 2590>
 "00000000000000000000101000011111", -- 2590 FREE #<CONS 0 2591>
 "00000000000000000000101000100000", -- 2591 FREE #<CONS 0 2592>
 "00000000000000000000101000100001", -- 2592 FREE #<CONS 0 2593>
 "00000000000000000000101000100010", -- 2593 FREE #<CONS 0 2594>
 "00000000000000000000101000100011", -- 2594 FREE #<CONS 0 2595>
 "00000000000000000000101000100100", -- 2595 FREE #<CONS 0 2596>
 "00000000000000000000101000100101", -- 2596 FREE #<CONS 0 2597>
 "00000000000000000000101000100110", -- 2597 FREE #<CONS 0 2598>
 "00000000000000000000101000100111", -- 2598 FREE #<CONS 0 2599>
 "00000000000000000000101000101000", -- 2599 FREE #<CONS 0 2600>
 "00000000000000000000101000101001", -- 2600 FREE #<CONS 0 2601>
 "00000000000000000000101000101010", -- 2601 FREE #<CONS 0 2602>
 "00000000000000000000101000101011", -- 2602 FREE #<CONS 0 2603>
 "00000000000000000000101000101100", -- 2603 FREE #<CONS 0 2604>
 "00000000000000000000101000101101", -- 2604 FREE #<CONS 0 2605>
 "00000000000000000000101000101110", -- 2605 FREE #<CONS 0 2606>
 "00000000000000000000101000101111", -- 2606 FREE #<CONS 0 2607>
 "00000000000000000000101000110000", -- 2607 FREE #<CONS 0 2608>
 "00000000000000000000101000110001", -- 2608 FREE #<CONS 0 2609>
 "00000000000000000000101000110010", -- 2609 FREE #<CONS 0 2610>
 "00000000000000000000101000110011", -- 2610 FREE #<CONS 0 2611>
 "00000000000000000000101000110100", -- 2611 FREE #<CONS 0 2612>
 "00000000000000000000101000110101", -- 2612 FREE #<CONS 0 2613>
 "00000000000000000000101000110110", -- 2613 FREE #<CONS 0 2614>
 "00000000000000000000101000110111", -- 2614 FREE #<CONS 0 2615>
 "00000000000000000000101000111000", -- 2615 FREE #<CONS 0 2616>
 "00000000000000000000101000111001", -- 2616 FREE #<CONS 0 2617>
 "00000000000000000000101000111010", -- 2617 FREE #<CONS 0 2618>
 "00000000000000000000101000111011", -- 2618 FREE #<CONS 0 2619>
 "00000000000000000000101000111100", -- 2619 FREE #<CONS 0 2620>
 "00000000000000000000101000111101", -- 2620 FREE #<CONS 0 2621>
 "00000000000000000000101000111110", -- 2621 FREE #<CONS 0 2622>
 "00000000000000000000101000111111", -- 2622 FREE #<CONS 0 2623>
 "00000000000000000000101001000000", -- 2623 FREE #<CONS 0 2624>
 "00000000000000000000101001000001", -- 2624 FREE #<CONS 0 2625>
 "00000000000000000000101001000010", -- 2625 FREE #<CONS 0 2626>
 "00000000000000000000101001000011", -- 2626 FREE #<CONS 0 2627>
 "00000000000000000000101001000100", -- 2627 FREE #<CONS 0 2628>
 "00000000000000000000101001000101", -- 2628 FREE #<CONS 0 2629>
 "00000000000000000000101001000110", -- 2629 FREE #<CONS 0 2630>
 "00000000000000000000101001000111", -- 2630 FREE #<CONS 0 2631>
 "00000000000000000000101001001000", -- 2631 FREE #<CONS 0 2632>
 "00000000000000000000101001001001", -- 2632 FREE #<CONS 0 2633>
 "00000000000000000000101001001010", -- 2633 FREE #<CONS 0 2634>
 "00000000000000000000101001001011", -- 2634 FREE #<CONS 0 2635>
 "00000000000000000000101001001100", -- 2635 FREE #<CONS 0 2636>
 "00000000000000000000101001001101", -- 2636 FREE #<CONS 0 2637>
 "00000000000000000000101001001110", -- 2637 FREE #<CONS 0 2638>
 "00000000000000000000101001001111", -- 2638 FREE #<CONS 0 2639>
 "00000000000000000000101001010000", -- 2639 FREE #<CONS 0 2640>
 "00000000000000000000101001010001", -- 2640 FREE #<CONS 0 2641>
 "00000000000000000000101001010010", -- 2641 FREE #<CONS 0 2642>
 "00000000000000000000101001010011", -- 2642 FREE #<CONS 0 2643>
 "00000000000000000000101001010100", -- 2643 FREE #<CONS 0 2644>
 "00000000000000000000101001010101", -- 2644 FREE #<CONS 0 2645>
 "00000000000000000000101001010110", -- 2645 FREE #<CONS 0 2646>
 "00000000000000000000101001010111", -- 2646 FREE #<CONS 0 2647>
 "00000000000000000000101001011000", -- 2647 FREE #<CONS 0 2648>
 "00000000000000000000101001011001", -- 2648 FREE #<CONS 0 2649>
 "00000000000000000000101001011010", -- 2649 FREE #<CONS 0 2650>
 "00000000000000000000101001011011", -- 2650 FREE #<CONS 0 2651>
 "00000000000000000000101001011100", -- 2651 FREE #<CONS 0 2652>
 "00000000000000000000101001011101", -- 2652 FREE #<CONS 0 2653>
 "00000000000000000000101001011110", -- 2653 FREE #<CONS 0 2654>
 "00000000000000000000101001011111", -- 2654 FREE #<CONS 0 2655>
 "00000000000000000000101001100000", -- 2655 FREE #<CONS 0 2656>
 "00000000000000000000101001100001", -- 2656 FREE #<CONS 0 2657>
 "00000000000000000000101001100010", -- 2657 FREE #<CONS 0 2658>
 "00000000000000000000101001100011", -- 2658 FREE #<CONS 0 2659>
 "00000000000000000000101001100100", -- 2659 FREE #<CONS 0 2660>
 "00000000000000000000101001100101", -- 2660 FREE #<CONS 0 2661>
 "00000000000000000000101001100110", -- 2661 FREE #<CONS 0 2662>
 "00000000000000000000101001100111", -- 2662 FREE #<CONS 0 2663>
 "00000000000000000000101001101000", -- 2663 FREE #<CONS 0 2664>
 "00000000000000000000101001101001", -- 2664 FREE #<CONS 0 2665>
 "00000000000000000000101001101010", -- 2665 FREE #<CONS 0 2666>
 "00000000000000000000101001101011", -- 2666 FREE #<CONS 0 2667>
 "00000000000000000000101001101100", -- 2667 FREE #<CONS 0 2668>
 "00000000000000000000101001101101", -- 2668 FREE #<CONS 0 2669>
 "00000000000000000000101001101110", -- 2669 FREE #<CONS 0 2670>
 "00000000000000000000101001101111", -- 2670 FREE #<CONS 0 2671>
 "00000000000000000000101001110000", -- 2671 FREE #<CONS 0 2672>
 "00000000000000000000101001110001", -- 2672 FREE #<CONS 0 2673>
 "00000000000000000000101001110010", -- 2673 FREE #<CONS 0 2674>
 "00000000000000000000101001110011", -- 2674 FREE #<CONS 0 2675>
 "00000000000000000000101001110100", -- 2675 FREE #<CONS 0 2676>
 "00000000000000000000101001110101", -- 2676 FREE #<CONS 0 2677>
 "00000000000000000000101001110110", -- 2677 FREE #<CONS 0 2678>
 "00000000000000000000101001110111", -- 2678 FREE #<CONS 0 2679>
 "00000000000000000000101001111000", -- 2679 FREE #<CONS 0 2680>
 "00000000000000000000101001111001", -- 2680 FREE #<CONS 0 2681>
 "00000000000000000000101001111010", -- 2681 FREE #<CONS 0 2682>
 "00000000000000000000101001111011", -- 2682 FREE #<CONS 0 2683>
 "00000000000000000000101001111100", -- 2683 FREE #<CONS 0 2684>
 "00000000000000000000101001111101", -- 2684 FREE #<CONS 0 2685>
 "00000000000000000000101001111110", -- 2685 FREE #<CONS 0 2686>
 "00000000000000000000101001111111", -- 2686 FREE #<CONS 0 2687>
 "00000000000000000000101010000000", -- 2687 FREE #<CONS 0 2688>
 "00000000000000000000101010000001", -- 2688 FREE #<CONS 0 2689>
 "00000000000000000000101010000010", -- 2689 FREE #<CONS 0 2690>
 "00000000000000000000101010000011", -- 2690 FREE #<CONS 0 2691>
 "00000000000000000000101010000100", -- 2691 FREE #<CONS 0 2692>
 "00000000000000000000101010000101", -- 2692 FREE #<CONS 0 2693>
 "00000000000000000000101010000110", -- 2693 FREE #<CONS 0 2694>
 "00000000000000000000101010000111", -- 2694 FREE #<CONS 0 2695>
 "00000000000000000000101010001000", -- 2695 FREE #<CONS 0 2696>
 "00000000000000000000101010001001", -- 2696 FREE #<CONS 0 2697>
 "00000000000000000000101010001010", -- 2697 FREE #<CONS 0 2698>
 "00000000000000000000101010001011", -- 2698 FREE #<CONS 0 2699>
 "00000000000000000000101010001100", -- 2699 FREE #<CONS 0 2700>
 "00000000000000000000101010001101", -- 2700 FREE #<CONS 0 2701>
 "00000000000000000000101010001110", -- 2701 FREE #<CONS 0 2702>
 "00000000000000000000101010001111", -- 2702 FREE #<CONS 0 2703>
 "00000000000000000000101010010000", -- 2703 FREE #<CONS 0 2704>
 "00000000000000000000101010010001", -- 2704 FREE #<CONS 0 2705>
 "00000000000000000000101010010010", -- 2705 FREE #<CONS 0 2706>
 "00000000000000000000101010010011", -- 2706 FREE #<CONS 0 2707>
 "00000000000000000000101010010100", -- 2707 FREE #<CONS 0 2708>
 "00000000000000000000101010010101", -- 2708 FREE #<CONS 0 2709>
 "00000000000000000000101010010110", -- 2709 FREE #<CONS 0 2710>
 "00000000000000000000101010010111", -- 2710 FREE #<CONS 0 2711>
 "00000000000000000000101010011000", -- 2711 FREE #<CONS 0 2712>
 "00000000000000000000101010011001", -- 2712 FREE #<CONS 0 2713>
 "00000000000000000000101010011010", -- 2713 FREE #<CONS 0 2714>
 "00000000000000000000101010011011", -- 2714 FREE #<CONS 0 2715>
 "00000000000000000000101010011100", -- 2715 FREE #<CONS 0 2716>
 "00000000000000000000101010011101", -- 2716 FREE #<CONS 0 2717>
 "00000000000000000000101010011110", -- 2717 FREE #<CONS 0 2718>
 "00000000000000000000101010011111", -- 2718 FREE #<CONS 0 2719>
 "00000000000000000000101010100000", -- 2719 FREE #<CONS 0 2720>
 "00000000000000000000101010100001", -- 2720 FREE #<CONS 0 2721>
 "00000000000000000000101010100010", -- 2721 FREE #<CONS 0 2722>
 "00000000000000000000101010100011", -- 2722 FREE #<CONS 0 2723>
 "00000000000000000000101010100100", -- 2723 FREE #<CONS 0 2724>
 "00000000000000000000101010100101", -- 2724 FREE #<CONS 0 2725>
 "00000000000000000000101010100110", -- 2725 FREE #<CONS 0 2726>
 "00000000000000000000101010100111", -- 2726 FREE #<CONS 0 2727>
 "00000000000000000000101010101000", -- 2727 FREE #<CONS 0 2728>
 "00000000000000000000101010101001", -- 2728 FREE #<CONS 0 2729>
 "00000000000000000000101010101010", -- 2729 FREE #<CONS 0 2730>
 "00000000000000000000101010101011", -- 2730 FREE #<CONS 0 2731>
 "00000000000000000000101010101100", -- 2731 FREE #<CONS 0 2732>
 "00000000000000000000101010101101", -- 2732 FREE #<CONS 0 2733>
 "00000000000000000000101010101110", -- 2733 FREE #<CONS 0 2734>
 "00000000000000000000101010101111", -- 2734 FREE #<CONS 0 2735>
 "00000000000000000000101010110000", -- 2735 FREE #<CONS 0 2736>
 "00000000000000000000101010110001", -- 2736 FREE #<CONS 0 2737>
 "00000000000000000000101010110010", -- 2737 FREE #<CONS 0 2738>
 "00000000000000000000101010110011", -- 2738 FREE #<CONS 0 2739>
 "00000000000000000000101010110100", -- 2739 FREE #<CONS 0 2740>
 "00000000000000000000101010110101", -- 2740 FREE #<CONS 0 2741>
 "00000000000000000000101010110110", -- 2741 FREE #<CONS 0 2742>
 "00000000000000000000101010110111", -- 2742 FREE #<CONS 0 2743>
 "00000000000000000000101010111000", -- 2743 FREE #<CONS 0 2744>
 "00000000000000000000101010111001", -- 2744 FREE #<CONS 0 2745>
 "00000000000000000000101010111010", -- 2745 FREE #<CONS 0 2746>
 "00000000000000000000101010111011", -- 2746 FREE #<CONS 0 2747>
 "00000000000000000000101010111100", -- 2747 FREE #<CONS 0 2748>
 "00000000000000000000101010111101", -- 2748 FREE #<CONS 0 2749>
 "00000000000000000000101010111110", -- 2749 FREE #<CONS 0 2750>
 "00000000000000000000101010111111", -- 2750 FREE #<CONS 0 2751>
 "00000000000000000000101011000000", -- 2751 FREE #<CONS 0 2752>
 "00000000000000000000101011000001", -- 2752 FREE #<CONS 0 2753>
 "00000000000000000000101011000010", -- 2753 FREE #<CONS 0 2754>
 "00000000000000000000101011000011", -- 2754 FREE #<CONS 0 2755>
 "00000000000000000000101011000100", -- 2755 FREE #<CONS 0 2756>
 "00000000000000000000101011000101", -- 2756 FREE #<CONS 0 2757>
 "00000000000000000000101011000110", -- 2757 FREE #<CONS 0 2758>
 "00000000000000000000101011000111", -- 2758 FREE #<CONS 0 2759>
 "00000000000000000000101011001000", -- 2759 FREE #<CONS 0 2760>
 "00000000000000000000101011001001", -- 2760 FREE #<CONS 0 2761>
 "00000000000000000000101011001010", -- 2761 FREE #<CONS 0 2762>
 "00000000000000000000101011001011", -- 2762 FREE #<CONS 0 2763>
 "00000000000000000000101011001100", -- 2763 FREE #<CONS 0 2764>
 "00000000000000000000101011001101", -- 2764 FREE #<CONS 0 2765>
 "00000000000000000000101011001110", -- 2765 FREE #<CONS 0 2766>
 "00000000000000000000101011001111", -- 2766 FREE #<CONS 0 2767>
 "00000000000000000000101011010000", -- 2767 FREE #<CONS 0 2768>
 "00000000000000000000101011010001", -- 2768 FREE #<CONS 0 2769>
 "00000000000000000000101011010010", -- 2769 FREE #<CONS 0 2770>
 "00000000000000000000101011010011", -- 2770 FREE #<CONS 0 2771>
 "00000000000000000000101011010100", -- 2771 FREE #<CONS 0 2772>
 "00000000000000000000101011010101", -- 2772 FREE #<CONS 0 2773>
 "00000000000000000000101011010110", -- 2773 FREE #<CONS 0 2774>
 "00000000000000000000101011010111", -- 2774 FREE #<CONS 0 2775>
 "00000000000000000000101011011000", -- 2775 FREE #<CONS 0 2776>
 "00000000000000000000101011011001", -- 2776 FREE #<CONS 0 2777>
 "00000000000000000000101011011010", -- 2777 FREE #<CONS 0 2778>
 "00000000000000000000101011011011", -- 2778 FREE #<CONS 0 2779>
 "00000000000000000000101011011100", -- 2779 FREE #<CONS 0 2780>
 "00000000000000000000101011011101", -- 2780 FREE #<CONS 0 2781>
 "00000000000000000000101011011110", -- 2781 FREE #<CONS 0 2782>
 "00000000000000000000101011011111", -- 2782 FREE #<CONS 0 2783>
 "00000000000000000000101011100000", -- 2783 FREE #<CONS 0 2784>
 "00000000000000000000101011100001", -- 2784 FREE #<CONS 0 2785>
 "00000000000000000000101011100010", -- 2785 FREE #<CONS 0 2786>
 "00000000000000000000101011100011", -- 2786 FREE #<CONS 0 2787>
 "00000000000000000000101011100100", -- 2787 FREE #<CONS 0 2788>
 "00000000000000000000101011100101", -- 2788 FREE #<CONS 0 2789>
 "00000000000000000000101011100110", -- 2789 FREE #<CONS 0 2790>
 "00000000000000000000101011100111", -- 2790 FREE #<CONS 0 2791>
 "00000000000000000000101011101000", -- 2791 FREE #<CONS 0 2792>
 "00000000000000000000101011101001", -- 2792 FREE #<CONS 0 2793>
 "00000000000000000000101011101010", -- 2793 FREE #<CONS 0 2794>
 "00000000000000000000101011101011", -- 2794 FREE #<CONS 0 2795>
 "00000000000000000000101011101100", -- 2795 FREE #<CONS 0 2796>
 "00000000000000000000101011101101", -- 2796 FREE #<CONS 0 2797>
 "00000000000000000000101011101110", -- 2797 FREE #<CONS 0 2798>
 "00000000000000000000101011101111", -- 2798 FREE #<CONS 0 2799>
 "00000000000000000000101011110000", -- 2799 FREE #<CONS 0 2800>
 "00000000000000000000101011110001", -- 2800 FREE #<CONS 0 2801>
 "00000000000000000000101011110010", -- 2801 FREE #<CONS 0 2802>
 "00000000000000000000101011110011", -- 2802 FREE #<CONS 0 2803>
 "00000000000000000000101011110100", -- 2803 FREE #<CONS 0 2804>
 "00000000000000000000101011110101", -- 2804 FREE #<CONS 0 2805>
 "00000000000000000000101011110110", -- 2805 FREE #<CONS 0 2806>
 "00000000000000000000101011110111", -- 2806 FREE #<CONS 0 2807>
 "00000000000000000000101011111000", -- 2807 FREE #<CONS 0 2808>
 "00000000000000000000101011111001", -- 2808 FREE #<CONS 0 2809>
 "00000000000000000000101011111010", -- 2809 FREE #<CONS 0 2810>
 "00000000000000000000101011111011", -- 2810 FREE #<CONS 0 2811>
 "00000000000000000000101011111100", -- 2811 FREE #<CONS 0 2812>
 "00000000000000000000101011111101", -- 2812 FREE #<CONS 0 2813>
 "00000000000000000000101011111110", -- 2813 FREE #<CONS 0 2814>
 "00000000000000000000101011111111", -- 2814 FREE #<CONS 0 2815>
 "00000000000000000000101100000000", -- 2815 FREE #<CONS 0 2816>
 "00000000000000000000101100000001", -- 2816 FREE #<CONS 0 2817>
 "00000000000000000000101100000010", -- 2817 FREE #<CONS 0 2818>
 "00000000000000000000101100000011", -- 2818 FREE #<CONS 0 2819>
 "00000000000000000000101100000100", -- 2819 FREE #<CONS 0 2820>
 "00000000000000000000101100000101", -- 2820 FREE #<CONS 0 2821>
 "00000000000000000000101100000110", -- 2821 FREE #<CONS 0 2822>
 "00000000000000000000101100000111", -- 2822 FREE #<CONS 0 2823>
 "00000000000000000000101100001000", -- 2823 FREE #<CONS 0 2824>
 "00000000000000000000101100001001", -- 2824 FREE #<CONS 0 2825>
 "00000000000000000000101100001010", -- 2825 FREE #<CONS 0 2826>
 "00000000000000000000101100001011", -- 2826 FREE #<CONS 0 2827>
 "00000000000000000000101100001100", -- 2827 FREE #<CONS 0 2828>
 "00000000000000000000101100001101", -- 2828 FREE #<CONS 0 2829>
 "00000000000000000000101100001110", -- 2829 FREE #<CONS 0 2830>
 "00000000000000000000101100001111", -- 2830 FREE #<CONS 0 2831>
 "00000000000000000000101100010000", -- 2831 FREE #<CONS 0 2832>
 "00000000000000000000101100010001", -- 2832 FREE #<CONS 0 2833>
 "00000000000000000000101100010010", -- 2833 FREE #<CONS 0 2834>
 "00000000000000000000101100010011", -- 2834 FREE #<CONS 0 2835>
 "00000000000000000000101100010100", -- 2835 FREE #<CONS 0 2836>
 "00000000000000000000101100010101", -- 2836 FREE #<CONS 0 2837>
 "00000000000000000000101100010110", -- 2837 FREE #<CONS 0 2838>
 "00000000000000000000101100010111", -- 2838 FREE #<CONS 0 2839>
 "00000000000000000000101100011000", -- 2839 FREE #<CONS 0 2840>
 "00000000000000000000101100011001", -- 2840 FREE #<CONS 0 2841>
 "00000000000000000000101100011010", -- 2841 FREE #<CONS 0 2842>
 "00000000000000000000101100011011", -- 2842 FREE #<CONS 0 2843>
 "00000000000000000000101100011100", -- 2843 FREE #<CONS 0 2844>
 "00000000000000000000101100011101", -- 2844 FREE #<CONS 0 2845>
 "00000000000000000000101100011110", -- 2845 FREE #<CONS 0 2846>
 "00000000000000000000101100011111", -- 2846 FREE #<CONS 0 2847>
 "00000000000000000000101100100000", -- 2847 FREE #<CONS 0 2848>
 "00000000000000000000101100100001", -- 2848 FREE #<CONS 0 2849>
 "00000000000000000000101100100010", -- 2849 FREE #<CONS 0 2850>
 "00000000000000000000101100100011", -- 2850 FREE #<CONS 0 2851>
 "00000000000000000000101100100100", -- 2851 FREE #<CONS 0 2852>
 "00000000000000000000101100100101", -- 2852 FREE #<CONS 0 2853>
 "00000000000000000000101100100110", -- 2853 FREE #<CONS 0 2854>
 "00000000000000000000101100100111", -- 2854 FREE #<CONS 0 2855>
 "00000000000000000000101100101000", -- 2855 FREE #<CONS 0 2856>
 "00000000000000000000101100101001", -- 2856 FREE #<CONS 0 2857>
 "00000000000000000000101100101010", -- 2857 FREE #<CONS 0 2858>
 "00000000000000000000101100101011", -- 2858 FREE #<CONS 0 2859>
 "00000000000000000000101100101100", -- 2859 FREE #<CONS 0 2860>
 "00000000000000000000101100101101", -- 2860 FREE #<CONS 0 2861>
 "00000000000000000000101100101110", -- 2861 FREE #<CONS 0 2862>
 "00000000000000000000101100101111", -- 2862 FREE #<CONS 0 2863>
 "00000000000000000000101100110000", -- 2863 FREE #<CONS 0 2864>
 "00000000000000000000101100110001", -- 2864 FREE #<CONS 0 2865>
 "00000000000000000000101100110010", -- 2865 FREE #<CONS 0 2866>
 "00000000000000000000101100110011", -- 2866 FREE #<CONS 0 2867>
 "00000000000000000000101100110100", -- 2867 FREE #<CONS 0 2868>
 "00000000000000000000101100110101", -- 2868 FREE #<CONS 0 2869>
 "00000000000000000000101100110110", -- 2869 FREE #<CONS 0 2870>
 "00000000000000000000101100110111", -- 2870 FREE #<CONS 0 2871>
 "00000000000000000000101100111000", -- 2871 FREE #<CONS 0 2872>
 "00000000000000000000101100111001", -- 2872 FREE #<CONS 0 2873>
 "00000000000000000000101100111010", -- 2873 FREE #<CONS 0 2874>
 "00000000000000000000101100111011", -- 2874 FREE #<CONS 0 2875>
 "00000000000000000000101100111100", -- 2875 FREE #<CONS 0 2876>
 "00000000000000000000101100111101", -- 2876 FREE #<CONS 0 2877>
 "00000000000000000000101100111110", -- 2877 FREE #<CONS 0 2878>
 "00000000000000000000101100111111", -- 2878 FREE #<CONS 0 2879>
 "00000000000000000000101101000000", -- 2879 FREE #<CONS 0 2880>
 "00000000000000000000101101000001", -- 2880 FREE #<CONS 0 2881>
 "00000000000000000000101101000010", -- 2881 FREE #<CONS 0 2882>
 "00000000000000000000101101000011", -- 2882 FREE #<CONS 0 2883>
 "00000000000000000000101101000100", -- 2883 FREE #<CONS 0 2884>
 "00000000000000000000101101000101", -- 2884 FREE #<CONS 0 2885>
 "00000000000000000000101101000110", -- 2885 FREE #<CONS 0 2886>
 "00000000000000000000101101000111", -- 2886 FREE #<CONS 0 2887>
 "00000000000000000000101101001000", -- 2887 FREE #<CONS 0 2888>
 "00000000000000000000101101001001", -- 2888 FREE #<CONS 0 2889>
 "00000000000000000000101101001010", -- 2889 FREE #<CONS 0 2890>
 "00000000000000000000101101001011", -- 2890 FREE #<CONS 0 2891>
 "00000000000000000000101101001100", -- 2891 FREE #<CONS 0 2892>
 "00000000000000000000101101001101", -- 2892 FREE #<CONS 0 2893>
 "00000000000000000000101101001110", -- 2893 FREE #<CONS 0 2894>
 "00000000000000000000101101001111", -- 2894 FREE #<CONS 0 2895>
 "00000000000000000000101101010000", -- 2895 FREE #<CONS 0 2896>
 "00000000000000000000101101010001", -- 2896 FREE #<CONS 0 2897>
 "00000000000000000000101101010010", -- 2897 FREE #<CONS 0 2898>
 "00000000000000000000101101010011", -- 2898 FREE #<CONS 0 2899>
 "00000000000000000000101101010100", -- 2899 FREE #<CONS 0 2900>
 "00000000000000000000101101010101", -- 2900 FREE #<CONS 0 2901>
 "00000000000000000000101101010110", -- 2901 FREE #<CONS 0 2902>
 "00000000000000000000101101010111", -- 2902 FREE #<CONS 0 2903>
 "00000000000000000000101101011000", -- 2903 FREE #<CONS 0 2904>
 "00000000000000000000101101011001", -- 2904 FREE #<CONS 0 2905>
 "00000000000000000000101101011010", -- 2905 FREE #<CONS 0 2906>
 "00000000000000000000101101011011", -- 2906 FREE #<CONS 0 2907>
 "00000000000000000000101101011100", -- 2907 FREE #<CONS 0 2908>
 "00000000000000000000101101011101", -- 2908 FREE #<CONS 0 2909>
 "00000000000000000000101101011110", -- 2909 FREE #<CONS 0 2910>
 "00000000000000000000101101011111", -- 2910 FREE #<CONS 0 2911>
 "00000000000000000000101101100000", -- 2911 FREE #<CONS 0 2912>
 "00000000000000000000101101100001", -- 2912 FREE #<CONS 0 2913>
 "00000000000000000000101101100010", -- 2913 FREE #<CONS 0 2914>
 "00000000000000000000101101100011", -- 2914 FREE #<CONS 0 2915>
 "00000000000000000000101101100100", -- 2915 FREE #<CONS 0 2916>
 "00000000000000000000101101100101", -- 2916 FREE #<CONS 0 2917>
 "00000000000000000000101101100110", -- 2917 FREE #<CONS 0 2918>
 "00000000000000000000101101100111", -- 2918 FREE #<CONS 0 2919>
 "00000000000000000000101101101000", -- 2919 FREE #<CONS 0 2920>
 "00000000000000000000101101101001", -- 2920 FREE #<CONS 0 2921>
 "00000000000000000000101101101010", -- 2921 FREE #<CONS 0 2922>
 "00000000000000000000101101101011", -- 2922 FREE #<CONS 0 2923>
 "00000000000000000000101101101100", -- 2923 FREE #<CONS 0 2924>
 "00000000000000000000101101101101", -- 2924 FREE #<CONS 0 2925>
 "00000000000000000000101101101110", -- 2925 FREE #<CONS 0 2926>
 "00000000000000000000101101101111", -- 2926 FREE #<CONS 0 2927>
 "00000000000000000000101101110000", -- 2927 FREE #<CONS 0 2928>
 "00000000000000000000101101110001", -- 2928 FREE #<CONS 0 2929>
 "00000000000000000000101101110010", -- 2929 FREE #<CONS 0 2930>
 "00000000000000000000101101110011", -- 2930 FREE #<CONS 0 2931>
 "00000000000000000000101101110100", -- 2931 FREE #<CONS 0 2932>
 "00000000000000000000101101110101", -- 2932 FREE #<CONS 0 2933>
 "00000000000000000000101101110110", -- 2933 FREE #<CONS 0 2934>
 "00000000000000000000101101110111", -- 2934 FREE #<CONS 0 2935>
 "00000000000000000000101101111000", -- 2935 FREE #<CONS 0 2936>
 "00000000000000000000101101111001", -- 2936 FREE #<CONS 0 2937>
 "00000000000000000000101101111010", -- 2937 FREE #<CONS 0 2938>
 "00000000000000000000101101111011", -- 2938 FREE #<CONS 0 2939>
 "00000000000000000000101101111100", -- 2939 FREE #<CONS 0 2940>
 "00000000000000000000101101111101", -- 2940 FREE #<CONS 0 2941>
 "00000000000000000000101101111110", -- 2941 FREE #<CONS 0 2942>
 "00000000000000000000101101111111", -- 2942 FREE #<CONS 0 2943>
 "00000000000000000000101110000000", -- 2943 FREE #<CONS 0 2944>
 "00000000000000000000101110000001", -- 2944 FREE #<CONS 0 2945>
 "00000000000000000000101110000010", -- 2945 FREE #<CONS 0 2946>
 "00000000000000000000101110000011", -- 2946 FREE #<CONS 0 2947>
 "00000000000000000000101110000100", -- 2947 FREE #<CONS 0 2948>
 "00000000000000000000101110000101", -- 2948 FREE #<CONS 0 2949>
 "00000000000000000000101110000110", -- 2949 FREE #<CONS 0 2950>
 "00000000000000000000101110000111", -- 2950 FREE #<CONS 0 2951>
 "00000000000000000000101110001000", -- 2951 FREE #<CONS 0 2952>
 "00000000000000000000101110001001", -- 2952 FREE #<CONS 0 2953>
 "00000000000000000000101110001010", -- 2953 FREE #<CONS 0 2954>
 "00000000000000000000101110001011", -- 2954 FREE #<CONS 0 2955>
 "00000000000000000000101110001100", -- 2955 FREE #<CONS 0 2956>
 "00000000000000000000101110001101", -- 2956 FREE #<CONS 0 2957>
 "00000000000000000000101110001110", -- 2957 FREE #<CONS 0 2958>
 "00000000000000000000101110001111", -- 2958 FREE #<CONS 0 2959>
 "00000000000000000000101110010000", -- 2959 FREE #<CONS 0 2960>
 "00000000000000000000101110010001", -- 2960 FREE #<CONS 0 2961>
 "00000000000000000000101110010010", -- 2961 FREE #<CONS 0 2962>
 "00000000000000000000101110010011", -- 2962 FREE #<CONS 0 2963>
 "00000000000000000000101110010100", -- 2963 FREE #<CONS 0 2964>
 "00000000000000000000101110010101", -- 2964 FREE #<CONS 0 2965>
 "00000000000000000000101110010110", -- 2965 FREE #<CONS 0 2966>
 "00000000000000000000101110010111", -- 2966 FREE #<CONS 0 2967>
 "00000000000000000000101110011000", -- 2967 FREE #<CONS 0 2968>
 "00000000000000000000101110011001", -- 2968 FREE #<CONS 0 2969>
 "00000000000000000000101110011010", -- 2969 FREE #<CONS 0 2970>
 "00000000000000000000101110011011", -- 2970 FREE #<CONS 0 2971>
 "00000000000000000000101110011100", -- 2971 FREE #<CONS 0 2972>
 "00000000000000000000101110011101", -- 2972 FREE #<CONS 0 2973>
 "00000000000000000000101110011110", -- 2973 FREE #<CONS 0 2974>
 "00000000000000000000101110011111", -- 2974 FREE #<CONS 0 2975>
 "00000000000000000000101110100000", -- 2975 FREE #<CONS 0 2976>
 "00000000000000000000101110100001", -- 2976 FREE #<CONS 0 2977>
 "00000000000000000000101110100010", -- 2977 FREE #<CONS 0 2978>
 "00000000000000000000101110100011", -- 2978 FREE #<CONS 0 2979>
 "00000000000000000000101110100100", -- 2979 FREE #<CONS 0 2980>
 "00000000000000000000101110100101", -- 2980 FREE #<CONS 0 2981>
 "00000000000000000000101110100110", -- 2981 FREE #<CONS 0 2982>
 "00000000000000000000101110100111", -- 2982 FREE #<CONS 0 2983>
 "00000000000000000000101110101000", -- 2983 FREE #<CONS 0 2984>
 "00000000000000000000101110101001", -- 2984 FREE #<CONS 0 2985>
 "00000000000000000000101110101010", -- 2985 FREE #<CONS 0 2986>
 "00000000000000000000101110101011", -- 2986 FREE #<CONS 0 2987>
 "00000000000000000000101110101100", -- 2987 FREE #<CONS 0 2988>
 "00000000000000000000101110101101", -- 2988 FREE #<CONS 0 2989>
 "00000000000000000000101110101110", -- 2989 FREE #<CONS 0 2990>
 "00000000000000000000101110101111", -- 2990 FREE #<CONS 0 2991>
 "00000000000000000000101110110000", -- 2991 FREE #<CONS 0 2992>
 "00000000000000000000101110110001", -- 2992 FREE #<CONS 0 2993>
 "00000000000000000000101110110010", -- 2993 FREE #<CONS 0 2994>
 "00000000000000000000101110110011", -- 2994 FREE #<CONS 0 2995>
 "00000000000000000000101110110100", -- 2995 FREE #<CONS 0 2996>
 "00000000000000000000101110110101", -- 2996 FREE #<CONS 0 2997>
 "00000000000000000000101110110110", -- 2997 FREE #<CONS 0 2998>
 "00000000000000000000101110110111", -- 2998 FREE #<CONS 0 2999>
 "00000000000000000000101110111000", -- 2999 FREE #<CONS 0 3000>
 "00000000000000000000101110111001", -- 3000 FREE #<CONS 0 3001>
 "00000000000000000000101110111010", -- 3001 FREE #<CONS 0 3002>
 "00000000000000000000101110111011", -- 3002 FREE #<CONS 0 3003>
 "00000000000000000000101110111100", -- 3003 FREE #<CONS 0 3004>
 "00000000000000000000101110111101", -- 3004 FREE #<CONS 0 3005>
 "00000000000000000000101110111110", -- 3005 FREE #<CONS 0 3006>
 "00000000000000000000101110111111", -- 3006 FREE #<CONS 0 3007>
 "00000000000000000000101111000000", -- 3007 FREE #<CONS 0 3008>
 "00000000000000000000101111000001", -- 3008 FREE #<CONS 0 3009>
 "00000000000000000000101111000010", -- 3009 FREE #<CONS 0 3010>
 "00000000000000000000101111000011", -- 3010 FREE #<CONS 0 3011>
 "00000000000000000000101111000100", -- 3011 FREE #<CONS 0 3012>
 "00000000000000000000101111000101", -- 3012 FREE #<CONS 0 3013>
 "00000000000000000000101111000110", -- 3013 FREE #<CONS 0 3014>
 "00000000000000000000101111000111", -- 3014 FREE #<CONS 0 3015>
 "00000000000000000000101111001000", -- 3015 FREE #<CONS 0 3016>
 "00000000000000000000101111001001", -- 3016 FREE #<CONS 0 3017>
 "00000000000000000000101111001010", -- 3017 FREE #<CONS 0 3018>
 "00000000000000000000101111001011", -- 3018 FREE #<CONS 0 3019>
 "00000000000000000000101111001100", -- 3019 FREE #<CONS 0 3020>
 "00000000000000000000101111001101", -- 3020 FREE #<CONS 0 3021>
 "00000000000000000000101111001110", -- 3021 FREE #<CONS 0 3022>
 "00000000000000000000101111001111", -- 3022 FREE #<CONS 0 3023>
 "00000000000000000000101111010000", -- 3023 FREE #<CONS 0 3024>
 "00000000000000000000101111010001", -- 3024 FREE #<CONS 0 3025>
 "00000000000000000000101111010010", -- 3025 FREE #<CONS 0 3026>
 "00000000000000000000101111010011", -- 3026 FREE #<CONS 0 3027>
 "00000000000000000000101111010100", -- 3027 FREE #<CONS 0 3028>
 "00000000000000000000101111010101", -- 3028 FREE #<CONS 0 3029>
 "00000000000000000000101111010110", -- 3029 FREE #<CONS 0 3030>
 "00000000000000000000101111010111", -- 3030 FREE #<CONS 0 3031>
 "00000000000000000000101111011000", -- 3031 FREE #<CONS 0 3032>
 "00000000000000000000101111011001", -- 3032 FREE #<CONS 0 3033>
 "00000000000000000000101111011010", -- 3033 FREE #<CONS 0 3034>
 "00000000000000000000101111011011", -- 3034 FREE #<CONS 0 3035>
 "00000000000000000000101111011100", -- 3035 FREE #<CONS 0 3036>
 "00000000000000000000101111011101", -- 3036 FREE #<CONS 0 3037>
 "00000000000000000000101111011110", -- 3037 FREE #<CONS 0 3038>
 "00000000000000000000101111011111", -- 3038 FREE #<CONS 0 3039>
 "00000000000000000000101111100000", -- 3039 FREE #<CONS 0 3040>
 "00000000000000000000101111100001", -- 3040 FREE #<CONS 0 3041>
 "00000000000000000000101111100010", -- 3041 FREE #<CONS 0 3042>
 "00000000000000000000101111100011", -- 3042 FREE #<CONS 0 3043>
 "00000000000000000000101111100100", -- 3043 FREE #<CONS 0 3044>
 "00000000000000000000101111100101", -- 3044 FREE #<CONS 0 3045>
 "00000000000000000000101111100110", -- 3045 FREE #<CONS 0 3046>
 "00000000000000000000101111100111", -- 3046 FREE #<CONS 0 3047>
 "00000000000000000000101111101000", -- 3047 FREE #<CONS 0 3048>
 "00000000000000000000101111101001", -- 3048 FREE #<CONS 0 3049>
 "00000000000000000000101111101010", -- 3049 FREE #<CONS 0 3050>
 "00000000000000000000101111101011", -- 3050 FREE #<CONS 0 3051>
 "00000000000000000000101111101100", -- 3051 FREE #<CONS 0 3052>
 "00000000000000000000101111101101", -- 3052 FREE #<CONS 0 3053>
 "00000000000000000000101111101110", -- 3053 FREE #<CONS 0 3054>
 "00000000000000000000101111101111", -- 3054 FREE #<CONS 0 3055>
 "00000000000000000000101111110000", -- 3055 FREE #<CONS 0 3056>
 "00000000000000000000101111110001", -- 3056 FREE #<CONS 0 3057>
 "00000000000000000000101111110010", -- 3057 FREE #<CONS 0 3058>
 "00000000000000000000101111110011", -- 3058 FREE #<CONS 0 3059>
 "00000000000000000000101111110100", -- 3059 FREE #<CONS 0 3060>
 "00000000000000000000101111110101", -- 3060 FREE #<CONS 0 3061>
 "00000000000000000000101111110110", -- 3061 FREE #<CONS 0 3062>
 "00000000000000000000101111110111", -- 3062 FREE #<CONS 0 3063>
 "00000000000000000000101111111000", -- 3063 FREE #<CONS 0 3064>
 "00000000000000000000101111111001", -- 3064 FREE #<CONS 0 3065>
 "00000000000000000000101111111010", -- 3065 FREE #<CONS 0 3066>
 "00000000000000000000101111111011", -- 3066 FREE #<CONS 0 3067>
 "00000000000000000000101111111100", -- 3067 FREE #<CONS 0 3068>
 "00000000000000000000101111111101", -- 3068 FREE #<CONS 0 3069>
 "00000000000000000000101111111110", -- 3069 FREE #<CONS 0 3070>
 "00000000000000000000101111111111", -- 3070 FREE #<CONS 0 3071>
 "00000000000000000000110000000000", -- 3071 FREE #<CONS 0 3072>
 "00000000000000000000110000000001", -- 3072 FREE #<CONS 0 3073>
 "00000000000000000000110000000010", -- 3073 FREE #<CONS 0 3074>
 "00000000000000000000110000000011", -- 3074 FREE #<CONS 0 3075>
 "00000000000000000000110000000100", -- 3075 FREE #<CONS 0 3076>
 "00000000000000000000110000000101", -- 3076 FREE #<CONS 0 3077>
 "00000000000000000000110000000110", -- 3077 FREE #<CONS 0 3078>
 "00000000000000000000110000000111", -- 3078 FREE #<CONS 0 3079>
 "00000000000000000000110000001000", -- 3079 FREE #<CONS 0 3080>
 "00000000000000000000110000001001", -- 3080 FREE #<CONS 0 3081>
 "00000000000000000000110000001010", -- 3081 FREE #<CONS 0 3082>
 "00000000000000000000110000001011", -- 3082 FREE #<CONS 0 3083>
 "00000000000000000000110000001100", -- 3083 FREE #<CONS 0 3084>
 "00000000000000000000110000001101", -- 3084 FREE #<CONS 0 3085>
 "00000000000000000000110000001110", -- 3085 FREE #<CONS 0 3086>
 "00000000000000000000110000001111", -- 3086 FREE #<CONS 0 3087>
 "00000000000000000000110000010000", -- 3087 FREE #<CONS 0 3088>
 "00000000000000000000110000010001", -- 3088 FREE #<CONS 0 3089>
 "00000000000000000000110000010010", -- 3089 FREE #<CONS 0 3090>
 "00000000000000000000110000010011", -- 3090 FREE #<CONS 0 3091>
 "00000000000000000000110000010100", -- 3091 FREE #<CONS 0 3092>
 "00000000000000000000110000010101", -- 3092 FREE #<CONS 0 3093>
 "00000000000000000000110000010110", -- 3093 FREE #<CONS 0 3094>
 "00000000000000000000110000010111", -- 3094 FREE #<CONS 0 3095>
 "00000000000000000000110000011000", -- 3095 FREE #<CONS 0 3096>
 "00000000000000000000110000011001", -- 3096 FREE #<CONS 0 3097>
 "00000000000000000000110000011010", -- 3097 FREE #<CONS 0 3098>
 "00000000000000000000110000011011", -- 3098 FREE #<CONS 0 3099>
 "00000000000000000000110000011100", -- 3099 FREE #<CONS 0 3100>
 "00000000000000000000110000011101", -- 3100 FREE #<CONS 0 3101>
 "00000000000000000000110000011110", -- 3101 FREE #<CONS 0 3102>
 "00000000000000000000110000011111", -- 3102 FREE #<CONS 0 3103>
 "00000000000000000000110000100000", -- 3103 FREE #<CONS 0 3104>
 "00000000000000000000110000100001", -- 3104 FREE #<CONS 0 3105>
 "00000000000000000000110000100010", -- 3105 FREE #<CONS 0 3106>
 "00000000000000000000110000100011", -- 3106 FREE #<CONS 0 3107>
 "00000000000000000000110000100100", -- 3107 FREE #<CONS 0 3108>
 "00000000000000000000110000100101", -- 3108 FREE #<CONS 0 3109>
 "00000000000000000000110000100110", -- 3109 FREE #<CONS 0 3110>
 "00000000000000000000110000100111", -- 3110 FREE #<CONS 0 3111>
 "00000000000000000000110000101000", -- 3111 FREE #<CONS 0 3112>
 "00000000000000000000110000101001", -- 3112 FREE #<CONS 0 3113>
 "00000000000000000000110000101010", -- 3113 FREE #<CONS 0 3114>
 "00000000000000000000110000101011", -- 3114 FREE #<CONS 0 3115>
 "00000000000000000000110000101100", -- 3115 FREE #<CONS 0 3116>
 "00000000000000000000110000101101", -- 3116 FREE #<CONS 0 3117>
 "00000000000000000000110000101110", -- 3117 FREE #<CONS 0 3118>
 "00000000000000000000110000101111", -- 3118 FREE #<CONS 0 3119>
 "00000000000000000000110000110000", -- 3119 FREE #<CONS 0 3120>
 "00000000000000000000110000110001", -- 3120 FREE #<CONS 0 3121>
 "00000000000000000000110000110010", -- 3121 FREE #<CONS 0 3122>
 "00000000000000000000110000110011", -- 3122 FREE #<CONS 0 3123>
 "00000000000000000000110000110100", -- 3123 FREE #<CONS 0 3124>
 "00000000000000000000110000110101", -- 3124 FREE #<CONS 0 3125>
 "00000000000000000000110000110110", -- 3125 FREE #<CONS 0 3126>
 "00000000000000000000110000110111", -- 3126 FREE #<CONS 0 3127>
 "00000000000000000000110000111000", -- 3127 FREE #<CONS 0 3128>
 "00000000000000000000110000111001", -- 3128 FREE #<CONS 0 3129>
 "00000000000000000000110000111010", -- 3129 FREE #<CONS 0 3130>
 "00000000000000000000110000111011", -- 3130 FREE #<CONS 0 3131>
 "00000000000000000000110000111100", -- 3131 FREE #<CONS 0 3132>
 "00000000000000000000110000111101", -- 3132 FREE #<CONS 0 3133>
 "00000000000000000000110000111110", -- 3133 FREE #<CONS 0 3134>
 "00000000000000000000110000111111", -- 3134 FREE #<CONS 0 3135>
 "00000000000000000000110001000000", -- 3135 FREE #<CONS 0 3136>
 "00000000000000000000110001000001", -- 3136 FREE #<CONS 0 3137>
 "00000000000000000000110001000010", -- 3137 FREE #<CONS 0 3138>
 "00000000000000000000110001000011", -- 3138 FREE #<CONS 0 3139>
 "00000000000000000000110001000100", -- 3139 FREE #<CONS 0 3140>
 "00000000000000000000110001000101", -- 3140 FREE #<CONS 0 3141>
 "00000000000000000000110001000110", -- 3141 FREE #<CONS 0 3142>
 "00000000000000000000110001000111", -- 3142 FREE #<CONS 0 3143>
 "00000000000000000000110001001000", -- 3143 FREE #<CONS 0 3144>
 "00000000000000000000110001001001", -- 3144 FREE #<CONS 0 3145>
 "00000000000000000000110001001010", -- 3145 FREE #<CONS 0 3146>
 "00000000000000000000110001001011", -- 3146 FREE #<CONS 0 3147>
 "00000000000000000000110001001100", -- 3147 FREE #<CONS 0 3148>
 "00000000000000000000110001001101", -- 3148 FREE #<CONS 0 3149>
 "00000000000000000000110001001110", -- 3149 FREE #<CONS 0 3150>
 "00000000000000000000110001001111", -- 3150 FREE #<CONS 0 3151>
 "00000000000000000000110001010000", -- 3151 FREE #<CONS 0 3152>
 "00000000000000000000110001010001", -- 3152 FREE #<CONS 0 3153>
 "00000000000000000000110001010010", -- 3153 FREE #<CONS 0 3154>
 "00000000000000000000110001010011", -- 3154 FREE #<CONS 0 3155>
 "00000000000000000000110001010100", -- 3155 FREE #<CONS 0 3156>
 "00000000000000000000110001010101", -- 3156 FREE #<CONS 0 3157>
 "00000000000000000000110001010110", -- 3157 FREE #<CONS 0 3158>
 "00000000000000000000110001010111", -- 3158 FREE #<CONS 0 3159>
 "00000000000000000000110001011000", -- 3159 FREE #<CONS 0 3160>
 "00000000000000000000110001011001", -- 3160 FREE #<CONS 0 3161>
 "00000000000000000000110001011010", -- 3161 FREE #<CONS 0 3162>
 "00000000000000000000110001011011", -- 3162 FREE #<CONS 0 3163>
 "00000000000000000000110001011100", -- 3163 FREE #<CONS 0 3164>
 "00000000000000000000110001011101", -- 3164 FREE #<CONS 0 3165>
 "00000000000000000000110001011110", -- 3165 FREE #<CONS 0 3166>
 "00000000000000000000110001011111", -- 3166 FREE #<CONS 0 3167>
 "00000000000000000000110001100000", -- 3167 FREE #<CONS 0 3168>
 "00000000000000000000110001100001", -- 3168 FREE #<CONS 0 3169>
 "00000000000000000000110001100010", -- 3169 FREE #<CONS 0 3170>
 "00000000000000000000110001100011", -- 3170 FREE #<CONS 0 3171>
 "00000000000000000000110001100100", -- 3171 FREE #<CONS 0 3172>
 "00000000000000000000110001100101", -- 3172 FREE #<CONS 0 3173>
 "00000000000000000000110001100110", -- 3173 FREE #<CONS 0 3174>
 "00000000000000000000110001100111", -- 3174 FREE #<CONS 0 3175>
 "00000000000000000000110001101000", -- 3175 FREE #<CONS 0 3176>
 "00000000000000000000110001101001", -- 3176 FREE #<CONS 0 3177>
 "00000000000000000000110001101010", -- 3177 FREE #<CONS 0 3178>
 "00000000000000000000110001101011", -- 3178 FREE #<CONS 0 3179>
 "00000000000000000000110001101100", -- 3179 FREE #<CONS 0 3180>
 "00000000000000000000110001101101", -- 3180 FREE #<CONS 0 3181>
 "00000000000000000000110001101110", -- 3181 FREE #<CONS 0 3182>
 "00000000000000000000110001101111", -- 3182 FREE #<CONS 0 3183>
 "00000000000000000000110001110000", -- 3183 FREE #<CONS 0 3184>
 "00000000000000000000110001110001", -- 3184 FREE #<CONS 0 3185>
 "00000000000000000000110001110010", -- 3185 FREE #<CONS 0 3186>
 "00000000000000000000110001110011", -- 3186 FREE #<CONS 0 3187>
 "00000000000000000000110001110100", -- 3187 FREE #<CONS 0 3188>
 "00000000000000000000110001110101", -- 3188 FREE #<CONS 0 3189>
 "00000000000000000000110001110110", -- 3189 FREE #<CONS 0 3190>
 "00000000000000000000110001110111", -- 3190 FREE #<CONS 0 3191>
 "00000000000000000000110001111000", -- 3191 FREE #<CONS 0 3192>
 "00000000000000000000110001111001", -- 3192 FREE #<CONS 0 3193>
 "00000000000000000000110001111010", -- 3193 FREE #<CONS 0 3194>
 "00000000000000000000110001111011", -- 3194 FREE #<CONS 0 3195>
 "00000000000000000000110001111100", -- 3195 FREE #<CONS 0 3196>
 "00000000000000000000110001111101", -- 3196 FREE #<CONS 0 3197>
 "00000000000000000000110001111110", -- 3197 FREE #<CONS 0 3198>
 "00000000000000000000110001111111", -- 3198 FREE #<CONS 0 3199>
 "00000000000000000000110010000000", -- 3199 FREE #<CONS 0 3200>
 "00000000000000000000110010000001", -- 3200 FREE #<CONS 0 3201>
 "00000000000000000000110010000010", -- 3201 FREE #<CONS 0 3202>
 "00000000000000000000110010000011", -- 3202 FREE #<CONS 0 3203>
 "00000000000000000000110010000100", -- 3203 FREE #<CONS 0 3204>
 "00000000000000000000110010000101", -- 3204 FREE #<CONS 0 3205>
 "00000000000000000000110010000110", -- 3205 FREE #<CONS 0 3206>
 "00000000000000000000110010000111", -- 3206 FREE #<CONS 0 3207>
 "00000000000000000000110010001000", -- 3207 FREE #<CONS 0 3208>
 "00000000000000000000110010001001", -- 3208 FREE #<CONS 0 3209>
 "00000000000000000000110010001010", -- 3209 FREE #<CONS 0 3210>
 "00000000000000000000110010001011", -- 3210 FREE #<CONS 0 3211>
 "00000000000000000000110010001100", -- 3211 FREE #<CONS 0 3212>
 "00000000000000000000110010001101", -- 3212 FREE #<CONS 0 3213>
 "00000000000000000000110010001110", -- 3213 FREE #<CONS 0 3214>
 "00000000000000000000110010001111", -- 3214 FREE #<CONS 0 3215>
 "00000000000000000000110010010000", -- 3215 FREE #<CONS 0 3216>
 "00000000000000000000110010010001", -- 3216 FREE #<CONS 0 3217>
 "00000000000000000000110010010010", -- 3217 FREE #<CONS 0 3218>
 "00000000000000000000110010010011", -- 3218 FREE #<CONS 0 3219>
 "00000000000000000000110010010100", -- 3219 FREE #<CONS 0 3220>
 "00000000000000000000110010010101", -- 3220 FREE #<CONS 0 3221>
 "00000000000000000000110010010110", -- 3221 FREE #<CONS 0 3222>
 "00000000000000000000110010010111", -- 3222 FREE #<CONS 0 3223>
 "00000000000000000000110010011000", -- 3223 FREE #<CONS 0 3224>
 "00000000000000000000110010011001", -- 3224 FREE #<CONS 0 3225>
 "00000000000000000000110010011010", -- 3225 FREE #<CONS 0 3226>
 "00000000000000000000110010011011", -- 3226 FREE #<CONS 0 3227>
 "00000000000000000000110010011100", -- 3227 FREE #<CONS 0 3228>
 "00000000000000000000110010011101", -- 3228 FREE #<CONS 0 3229>
 "00000000000000000000110010011110", -- 3229 FREE #<CONS 0 3230>
 "00000000000000000000110010011111", -- 3230 FREE #<CONS 0 3231>
 "00000000000000000000110010100000", -- 3231 FREE #<CONS 0 3232>
 "00000000000000000000110010100001", -- 3232 FREE #<CONS 0 3233>
 "00000000000000000000110010100010", -- 3233 FREE #<CONS 0 3234>
 "00000000000000000000110010100011", -- 3234 FREE #<CONS 0 3235>
 "00000000000000000000110010100100", -- 3235 FREE #<CONS 0 3236>
 "00000000000000000000110010100101", -- 3236 FREE #<CONS 0 3237>
 "00000000000000000000110010100110", -- 3237 FREE #<CONS 0 3238>
 "00000000000000000000110010100111", -- 3238 FREE #<CONS 0 3239>
 "00000000000000000000110010101000", -- 3239 FREE #<CONS 0 3240>
 "00000000000000000000110010101001", -- 3240 FREE #<CONS 0 3241>
 "00000000000000000000110010101010", -- 3241 FREE #<CONS 0 3242>
 "00000000000000000000110010101011", -- 3242 FREE #<CONS 0 3243>
 "00000000000000000000110010101100", -- 3243 FREE #<CONS 0 3244>
 "00000000000000000000110010101101", -- 3244 FREE #<CONS 0 3245>
 "00000000000000000000110010101110", -- 3245 FREE #<CONS 0 3246>
 "00000000000000000000110010101111", -- 3246 FREE #<CONS 0 3247>
 "00000000000000000000110010110000", -- 3247 FREE #<CONS 0 3248>
 "00000000000000000000110010110001", -- 3248 FREE #<CONS 0 3249>
 "00000000000000000000110010110010", -- 3249 FREE #<CONS 0 3250>
 "00000000000000000000110010110011", -- 3250 FREE #<CONS 0 3251>
 "00000000000000000000110010110100", -- 3251 FREE #<CONS 0 3252>
 "00000000000000000000110010110101", -- 3252 FREE #<CONS 0 3253>
 "00000000000000000000110010110110", -- 3253 FREE #<CONS 0 3254>
 "00000000000000000000110010110111", -- 3254 FREE #<CONS 0 3255>
 "00000000000000000000110010111000", -- 3255 FREE #<CONS 0 3256>
 "00000000000000000000110010111001", -- 3256 FREE #<CONS 0 3257>
 "00000000000000000000110010111010", -- 3257 FREE #<CONS 0 3258>
 "00000000000000000000110010111011", -- 3258 FREE #<CONS 0 3259>
 "00000000000000000000110010111100", -- 3259 FREE #<CONS 0 3260>
 "00000000000000000000110010111101", -- 3260 FREE #<CONS 0 3261>
 "00000000000000000000110010111110", -- 3261 FREE #<CONS 0 3262>
 "00000000000000000000110010111111", -- 3262 FREE #<CONS 0 3263>
 "00000000000000000000110011000000", -- 3263 FREE #<CONS 0 3264>
 "00000000000000000000110011000001", -- 3264 FREE #<CONS 0 3265>
 "00000000000000000000110011000010", -- 3265 FREE #<CONS 0 3266>
 "00000000000000000000110011000011", -- 3266 FREE #<CONS 0 3267>
 "00000000000000000000110011000100", -- 3267 FREE #<CONS 0 3268>
 "00000000000000000000110011000101", -- 3268 FREE #<CONS 0 3269>
 "00000000000000000000110011000110", -- 3269 FREE #<CONS 0 3270>
 "00000000000000000000110011000111", -- 3270 FREE #<CONS 0 3271>
 "00000000000000000000110011001000", -- 3271 FREE #<CONS 0 3272>
 "00000000000000000000110011001001", -- 3272 FREE #<CONS 0 3273>
 "00000000000000000000110011001010", -- 3273 FREE #<CONS 0 3274>
 "00000000000000000000110011001011", -- 3274 FREE #<CONS 0 3275>
 "00000000000000000000110011001100", -- 3275 FREE #<CONS 0 3276>
 "00000000000000000000110011001101", -- 3276 FREE #<CONS 0 3277>
 "00000000000000000000110011001110", -- 3277 FREE #<CONS 0 3278>
 "00000000000000000000110011001111", -- 3278 FREE #<CONS 0 3279>
 "00000000000000000000110011010000", -- 3279 FREE #<CONS 0 3280>
 "00000000000000000000110011010001", -- 3280 FREE #<CONS 0 3281>
 "00000000000000000000110011010010", -- 3281 FREE #<CONS 0 3282>
 "00000000000000000000110011010011", -- 3282 FREE #<CONS 0 3283>
 "00000000000000000000110011010100", -- 3283 FREE #<CONS 0 3284>
 "00000000000000000000110011010101", -- 3284 FREE #<CONS 0 3285>
 "00000000000000000000110011010110", -- 3285 FREE #<CONS 0 3286>
 "00000000000000000000110011010111", -- 3286 FREE #<CONS 0 3287>
 "00000000000000000000110011011000", -- 3287 FREE #<CONS 0 3288>
 "00000000000000000000110011011001", -- 3288 FREE #<CONS 0 3289>
 "00000000000000000000110011011010", -- 3289 FREE #<CONS 0 3290>
 "00000000000000000000110011011011", -- 3290 FREE #<CONS 0 3291>
 "00000000000000000000110011011100", -- 3291 FREE #<CONS 0 3292>
 "00000000000000000000110011011101", -- 3292 FREE #<CONS 0 3293>
 "00000000000000000000110011011110", -- 3293 FREE #<CONS 0 3294>
 "00000000000000000000110011011111", -- 3294 FREE #<CONS 0 3295>
 "00000000000000000000110011100000", -- 3295 FREE #<CONS 0 3296>
 "00000000000000000000110011100001", -- 3296 FREE #<CONS 0 3297>
 "00000000000000000000110011100010", -- 3297 FREE #<CONS 0 3298>
 "00000000000000000000110011100011", -- 3298 FREE #<CONS 0 3299>
 "00000000000000000000110011100100", -- 3299 FREE #<CONS 0 3300>
 "00000000000000000000110011100101", -- 3300 FREE #<CONS 0 3301>
 "00000000000000000000110011100110", -- 3301 FREE #<CONS 0 3302>
 "00000000000000000000110011100111", -- 3302 FREE #<CONS 0 3303>
 "00000000000000000000110011101000", -- 3303 FREE #<CONS 0 3304>
 "00000000000000000000110011101001", -- 3304 FREE #<CONS 0 3305>
 "00000000000000000000110011101010", -- 3305 FREE #<CONS 0 3306>
 "00000000000000000000110011101011", -- 3306 FREE #<CONS 0 3307>
 "00000000000000000000110011101100", -- 3307 FREE #<CONS 0 3308>
 "00000000000000000000110011101101", -- 3308 FREE #<CONS 0 3309>
 "00000000000000000000110011101110", -- 3309 FREE #<CONS 0 3310>
 "00000000000000000000110011101111", -- 3310 FREE #<CONS 0 3311>
 "00000000000000000000110011110000", -- 3311 FREE #<CONS 0 3312>
 "00000000000000000000110011110001", -- 3312 FREE #<CONS 0 3313>
 "00000000000000000000110011110010", -- 3313 FREE #<CONS 0 3314>
 "00000000000000000000110011110011", -- 3314 FREE #<CONS 0 3315>
 "00000000000000000000110011110100", -- 3315 FREE #<CONS 0 3316>
 "00000000000000000000110011110101", -- 3316 FREE #<CONS 0 3317>
 "00000000000000000000110011110110", -- 3317 FREE #<CONS 0 3318>
 "00000000000000000000110011110111", -- 3318 FREE #<CONS 0 3319>
 "00000000000000000000110011111000", -- 3319 FREE #<CONS 0 3320>
 "00000000000000000000110011111001", -- 3320 FREE #<CONS 0 3321>
 "00000000000000000000110011111010", -- 3321 FREE #<CONS 0 3322>
 "00000000000000000000110011111011", -- 3322 FREE #<CONS 0 3323>
 "00000000000000000000110011111100", -- 3323 FREE #<CONS 0 3324>
 "00000000000000000000110011111101", -- 3324 FREE #<CONS 0 3325>
 "00000000000000000000110011111110", -- 3325 FREE #<CONS 0 3326>
 "00000000000000000000110011111111", -- 3326 FREE #<CONS 0 3327>
 "00000000000000000000110100000000", -- 3327 FREE #<CONS 0 3328>
 "00000000000000000000110100000001", -- 3328 FREE #<CONS 0 3329>
 "00000000000000000000110100000010", -- 3329 FREE #<CONS 0 3330>
 "00000000000000000000110100000011", -- 3330 FREE #<CONS 0 3331>
 "00000000000000000000110100000100", -- 3331 FREE #<CONS 0 3332>
 "00000000000000000000110100000101", -- 3332 FREE #<CONS 0 3333>
 "00000000000000000000110100000110", -- 3333 FREE #<CONS 0 3334>
 "00000000000000000000110100000111", -- 3334 FREE #<CONS 0 3335>
 "00000000000000000000110100001000", -- 3335 FREE #<CONS 0 3336>
 "00000000000000000000110100001001", -- 3336 FREE #<CONS 0 3337>
 "00000000000000000000110100001010", -- 3337 FREE #<CONS 0 3338>
 "00000000000000000000110100001011", -- 3338 FREE #<CONS 0 3339>
 "00000000000000000000110100001100", -- 3339 FREE #<CONS 0 3340>
 "00000000000000000000110100001101", -- 3340 FREE #<CONS 0 3341>
 "00000000000000000000110100001110", -- 3341 FREE #<CONS 0 3342>
 "00000000000000000000110100001111", -- 3342 FREE #<CONS 0 3343>
 "00000000000000000000110100010000", -- 3343 FREE #<CONS 0 3344>
 "00000000000000000000110100010001", -- 3344 FREE #<CONS 0 3345>
 "00000000000000000000110100010010", -- 3345 FREE #<CONS 0 3346>
 "00000000000000000000110100010011", -- 3346 FREE #<CONS 0 3347>
 "00000000000000000000110100010100", -- 3347 FREE #<CONS 0 3348>
 "00000000000000000000110100010101", -- 3348 FREE #<CONS 0 3349>
 "00000000000000000000110100010110", -- 3349 FREE #<CONS 0 3350>
 "00000000000000000000110100010111", -- 3350 FREE #<CONS 0 3351>
 "00000000000000000000110100011000", -- 3351 FREE #<CONS 0 3352>
 "00000000000000000000110100011001", -- 3352 FREE #<CONS 0 3353>
 "00000000000000000000110100011010", -- 3353 FREE #<CONS 0 3354>
 "00000000000000000000110100011011", -- 3354 FREE #<CONS 0 3355>
 "00000000000000000000110100011100", -- 3355 FREE #<CONS 0 3356>
 "00000000000000000000110100011101", -- 3356 FREE #<CONS 0 3357>
 "00000000000000000000110100011110", -- 3357 FREE #<CONS 0 3358>
 "00000000000000000000110100011111", -- 3358 FREE #<CONS 0 3359>
 "00000000000000000000110100100000", -- 3359 FREE #<CONS 0 3360>
 "00000000000000000000110100100001", -- 3360 FREE #<CONS 0 3361>
 "00000000000000000000110100100010", -- 3361 FREE #<CONS 0 3362>
 "00000000000000000000110100100011", -- 3362 FREE #<CONS 0 3363>
 "00000000000000000000110100100100", -- 3363 FREE #<CONS 0 3364>
 "00000000000000000000110100100101", -- 3364 FREE #<CONS 0 3365>
 "00000000000000000000110100100110", -- 3365 FREE #<CONS 0 3366>
 "00000000000000000000110100100111", -- 3366 FREE #<CONS 0 3367>
 "00000000000000000000110100101000", -- 3367 FREE #<CONS 0 3368>
 "00000000000000000000110100101001", -- 3368 FREE #<CONS 0 3369>
 "00000000000000000000110100101010", -- 3369 FREE #<CONS 0 3370>
 "00000000000000000000110100101011", -- 3370 FREE #<CONS 0 3371>
 "00000000000000000000110100101100", -- 3371 FREE #<CONS 0 3372>
 "00000000000000000000110100101101", -- 3372 FREE #<CONS 0 3373>
 "00000000000000000000110100101110", -- 3373 FREE #<CONS 0 3374>
 "00000000000000000000110100101111", -- 3374 FREE #<CONS 0 3375>
 "00000000000000000000110100110000", -- 3375 FREE #<CONS 0 3376>
 "00000000000000000000110100110001", -- 3376 FREE #<CONS 0 3377>
 "00000000000000000000110100110010", -- 3377 FREE #<CONS 0 3378>
 "00000000000000000000110100110011", -- 3378 FREE #<CONS 0 3379>
 "00000000000000000000110100110100", -- 3379 FREE #<CONS 0 3380>
 "00000000000000000000110100110101", -- 3380 FREE #<CONS 0 3381>
 "00000000000000000000110100110110", -- 3381 FREE #<CONS 0 3382>
 "00000000000000000000110100110111", -- 3382 FREE #<CONS 0 3383>
 "00000000000000000000110100111000", -- 3383 FREE #<CONS 0 3384>
 "00000000000000000000110100111001", -- 3384 FREE #<CONS 0 3385>
 "00000000000000000000110100111010", -- 3385 FREE #<CONS 0 3386>
 "00000000000000000000110100111011", -- 3386 FREE #<CONS 0 3387>
 "00000000000000000000110100111100", -- 3387 FREE #<CONS 0 3388>
 "00000000000000000000110100111101", -- 3388 FREE #<CONS 0 3389>
 "00000000000000000000110100111110", -- 3389 FREE #<CONS 0 3390>
 "00000000000000000000110100111111", -- 3390 FREE #<CONS 0 3391>
 "00000000000000000000110101000000", -- 3391 FREE #<CONS 0 3392>
 "00000000000000000000110101000001", -- 3392 FREE #<CONS 0 3393>
 "00000000000000000000110101000010", -- 3393 FREE #<CONS 0 3394>
 "00000000000000000000110101000011", -- 3394 FREE #<CONS 0 3395>
 "00000000000000000000110101000100", -- 3395 FREE #<CONS 0 3396>
 "00000000000000000000110101000101", -- 3396 FREE #<CONS 0 3397>
 "00000000000000000000110101000110", -- 3397 FREE #<CONS 0 3398>
 "00000000000000000000110101000111", -- 3398 FREE #<CONS 0 3399>
 "00000000000000000000110101001000", -- 3399 FREE #<CONS 0 3400>
 "00000000000000000000110101001001", -- 3400 FREE #<CONS 0 3401>
 "00000000000000000000110101001010", -- 3401 FREE #<CONS 0 3402>
 "00000000000000000000110101001011", -- 3402 FREE #<CONS 0 3403>
 "00000000000000000000110101001100", -- 3403 FREE #<CONS 0 3404>
 "00000000000000000000110101001101", -- 3404 FREE #<CONS 0 3405>
 "00000000000000000000110101001110", -- 3405 FREE #<CONS 0 3406>
 "00000000000000000000110101001111", -- 3406 FREE #<CONS 0 3407>
 "00000000000000000000110101010000", -- 3407 FREE #<CONS 0 3408>
 "00000000000000000000110101010001", -- 3408 FREE #<CONS 0 3409>
 "00000000000000000000110101010010", -- 3409 FREE #<CONS 0 3410>
 "00000000000000000000110101010011", -- 3410 FREE #<CONS 0 3411>
 "00000000000000000000110101010100", -- 3411 FREE #<CONS 0 3412>
 "00000000000000000000110101010101", -- 3412 FREE #<CONS 0 3413>
 "00000000000000000000110101010110", -- 3413 FREE #<CONS 0 3414>
 "00000000000000000000110101010111", -- 3414 FREE #<CONS 0 3415>
 "00000000000000000000110101011000", -- 3415 FREE #<CONS 0 3416>
 "00000000000000000000110101011001", -- 3416 FREE #<CONS 0 3417>
 "00000000000000000000110101011010", -- 3417 FREE #<CONS 0 3418>
 "00000000000000000000110101011011", -- 3418 FREE #<CONS 0 3419>
 "00000000000000000000110101011100", -- 3419 FREE #<CONS 0 3420>
 "00000000000000000000110101011101", -- 3420 FREE #<CONS 0 3421>
 "00000000000000000000110101011110", -- 3421 FREE #<CONS 0 3422>
 "00000000000000000000110101011111", -- 3422 FREE #<CONS 0 3423>
 "00000000000000000000110101100000", -- 3423 FREE #<CONS 0 3424>
 "00000000000000000000110101100001", -- 3424 FREE #<CONS 0 3425>
 "00000000000000000000110101100010", -- 3425 FREE #<CONS 0 3426>
 "00000000000000000000110101100011", -- 3426 FREE #<CONS 0 3427>
 "00000000000000000000110101100100", -- 3427 FREE #<CONS 0 3428>
 "00000000000000000000110101100101", -- 3428 FREE #<CONS 0 3429>
 "00000000000000000000110101100110", -- 3429 FREE #<CONS 0 3430>
 "00000000000000000000110101100111", -- 3430 FREE #<CONS 0 3431>
 "00000000000000000000110101101000", -- 3431 FREE #<CONS 0 3432>
 "00000000000000000000110101101001", -- 3432 FREE #<CONS 0 3433>
 "00000000000000000000110101101010", -- 3433 FREE #<CONS 0 3434>
 "00000000000000000000110101101011", -- 3434 FREE #<CONS 0 3435>
 "00000000000000000000110101101100", -- 3435 FREE #<CONS 0 3436>
 "00000000000000000000110101101101", -- 3436 FREE #<CONS 0 3437>
 "00000000000000000000110101101110", -- 3437 FREE #<CONS 0 3438>
 "00000000000000000000110101101111", -- 3438 FREE #<CONS 0 3439>
 "00000000000000000000110101110000", -- 3439 FREE #<CONS 0 3440>
 "00000000000000000000110101110001", -- 3440 FREE #<CONS 0 3441>
 "00000000000000000000110101110010", -- 3441 FREE #<CONS 0 3442>
 "00000000000000000000110101110011", -- 3442 FREE #<CONS 0 3443>
 "00000000000000000000110101110100", -- 3443 FREE #<CONS 0 3444>
 "00000000000000000000110101110101", -- 3444 FREE #<CONS 0 3445>
 "00000000000000000000110101110110", -- 3445 FREE #<CONS 0 3446>
 "00000000000000000000110101110111", -- 3446 FREE #<CONS 0 3447>
 "00000000000000000000110101111000", -- 3447 FREE #<CONS 0 3448>
 "00000000000000000000110101111001", -- 3448 FREE #<CONS 0 3449>
 "00000000000000000000110101111010", -- 3449 FREE #<CONS 0 3450>
 "00000000000000000000110101111011", -- 3450 FREE #<CONS 0 3451>
 "00000000000000000000110101111100", -- 3451 FREE #<CONS 0 3452>
 "00000000000000000000110101111101", -- 3452 FREE #<CONS 0 3453>
 "00000000000000000000110101111110", -- 3453 FREE #<CONS 0 3454>
 "00000000000000000000110101111111", -- 3454 FREE #<CONS 0 3455>
 "00000000000000000000110110000000", -- 3455 FREE #<CONS 0 3456>
 "00000000000000000000110110000001", -- 3456 FREE #<CONS 0 3457>
 "00000000000000000000110110000010", -- 3457 FREE #<CONS 0 3458>
 "00000000000000000000110110000011", -- 3458 FREE #<CONS 0 3459>
 "00000000000000000000110110000100", -- 3459 FREE #<CONS 0 3460>
 "00000000000000000000110110000101", -- 3460 FREE #<CONS 0 3461>
 "00000000000000000000110110000110", -- 3461 FREE #<CONS 0 3462>
 "00000000000000000000110110000111", -- 3462 FREE #<CONS 0 3463>
 "00000000000000000000110110001000", -- 3463 FREE #<CONS 0 3464>
 "00000000000000000000110110001001", -- 3464 FREE #<CONS 0 3465>
 "00000000000000000000110110001010", -- 3465 FREE #<CONS 0 3466>
 "00000000000000000000110110001011", -- 3466 FREE #<CONS 0 3467>
 "00000000000000000000110110001100", -- 3467 FREE #<CONS 0 3468>
 "00000000000000000000110110001101", -- 3468 FREE #<CONS 0 3469>
 "00000000000000000000110110001110", -- 3469 FREE #<CONS 0 3470>
 "00000000000000000000110110001111", -- 3470 FREE #<CONS 0 3471>
 "00000000000000000000110110010000", -- 3471 FREE #<CONS 0 3472>
 "00000000000000000000110110010001", -- 3472 FREE #<CONS 0 3473>
 "00000000000000000000110110010010", -- 3473 FREE #<CONS 0 3474>
 "00000000000000000000110110010011", -- 3474 FREE #<CONS 0 3475>
 "00000000000000000000110110010100", -- 3475 FREE #<CONS 0 3476>
 "00000000000000000000110110010101", -- 3476 FREE #<CONS 0 3477>
 "00000000000000000000110110010110", -- 3477 FREE #<CONS 0 3478>
 "00000000000000000000110110010111", -- 3478 FREE #<CONS 0 3479>
 "00000000000000000000110110011000", -- 3479 FREE #<CONS 0 3480>
 "00000000000000000000110110011001", -- 3480 FREE #<CONS 0 3481>
 "00000000000000000000110110011010", -- 3481 FREE #<CONS 0 3482>
 "00000000000000000000110110011011", -- 3482 FREE #<CONS 0 3483>
 "00000000000000000000110110011100", -- 3483 FREE #<CONS 0 3484>
 "00000000000000000000110110011101", -- 3484 FREE #<CONS 0 3485>
 "00000000000000000000110110011110", -- 3485 FREE #<CONS 0 3486>
 "00000000000000000000110110011111", -- 3486 FREE #<CONS 0 3487>
 "00000000000000000000110110100000", -- 3487 FREE #<CONS 0 3488>
 "00000000000000000000110110100001", -- 3488 FREE #<CONS 0 3489>
 "00000000000000000000110110100010", -- 3489 FREE #<CONS 0 3490>
 "00000000000000000000110110100011", -- 3490 FREE #<CONS 0 3491>
 "00000000000000000000110110100100", -- 3491 FREE #<CONS 0 3492>
 "00000000000000000000110110100101", -- 3492 FREE #<CONS 0 3493>
 "00000000000000000000110110100110", -- 3493 FREE #<CONS 0 3494>
 "00000000000000000000110110100111", -- 3494 FREE #<CONS 0 3495>
 "00000000000000000000110110101000", -- 3495 FREE #<CONS 0 3496>
 "00000000000000000000110110101001", -- 3496 FREE #<CONS 0 3497>
 "00000000000000000000110110101010", -- 3497 FREE #<CONS 0 3498>
 "00000000000000000000110110101011", -- 3498 FREE #<CONS 0 3499>
 "00000000000000000000110110101100", -- 3499 FREE #<CONS 0 3500>
 "00000000000000000000110110101101", -- 3500 FREE #<CONS 0 3501>
 "00000000000000000000110110101110", -- 3501 FREE #<CONS 0 3502>
 "00000000000000000000110110101111", -- 3502 FREE #<CONS 0 3503>
 "00000000000000000000110110110000", -- 3503 FREE #<CONS 0 3504>
 "00000000000000000000110110110001", -- 3504 FREE #<CONS 0 3505>
 "00000000000000000000110110110010", -- 3505 FREE #<CONS 0 3506>
 "00000000000000000000110110110011", -- 3506 FREE #<CONS 0 3507>
 "00000000000000000000110110110100", -- 3507 FREE #<CONS 0 3508>
 "00000000000000000000110110110101", -- 3508 FREE #<CONS 0 3509>
 "00000000000000000000110110110110", -- 3509 FREE #<CONS 0 3510>
 "00000000000000000000110110110111", -- 3510 FREE #<CONS 0 3511>
 "00000000000000000000110110111000", -- 3511 FREE #<CONS 0 3512>
 "00000000000000000000110110111001", -- 3512 FREE #<CONS 0 3513>
 "00000000000000000000110110111010", -- 3513 FREE #<CONS 0 3514>
 "00000000000000000000110110111011", -- 3514 FREE #<CONS 0 3515>
 "00000000000000000000110110111100", -- 3515 FREE #<CONS 0 3516>
 "00000000000000000000110110111101", -- 3516 FREE #<CONS 0 3517>
 "00000000000000000000110110111110", -- 3517 FREE #<CONS 0 3518>
 "00000000000000000000110110111111", -- 3518 FREE #<CONS 0 3519>
 "00000000000000000000110111000000", -- 3519 FREE #<CONS 0 3520>
 "00000000000000000000110111000001", -- 3520 FREE #<CONS 0 3521>
 "00000000000000000000110111000010", -- 3521 FREE #<CONS 0 3522>
 "00000000000000000000110111000011", -- 3522 FREE #<CONS 0 3523>
 "00000000000000000000110111000100", -- 3523 FREE #<CONS 0 3524>
 "00000000000000000000110111000101", -- 3524 FREE #<CONS 0 3525>
 "00000000000000000000110111000110", -- 3525 FREE #<CONS 0 3526>
 "00000000000000000000110111000111", -- 3526 FREE #<CONS 0 3527>
 "00000000000000000000110111001000", -- 3527 FREE #<CONS 0 3528>
 "00000000000000000000110111001001", -- 3528 FREE #<CONS 0 3529>
 "00000000000000000000110111001010", -- 3529 FREE #<CONS 0 3530>
 "00000000000000000000110111001011", -- 3530 FREE #<CONS 0 3531>
 "00000000000000000000110111001100", -- 3531 FREE #<CONS 0 3532>
 "00000000000000000000110111001101", -- 3532 FREE #<CONS 0 3533>
 "00000000000000000000110111001110", -- 3533 FREE #<CONS 0 3534>
 "00000000000000000000110111001111", -- 3534 FREE #<CONS 0 3535>
 "00000000000000000000110111010000", -- 3535 FREE #<CONS 0 3536>
 "00000000000000000000110111010001", -- 3536 FREE #<CONS 0 3537>
 "00000000000000000000110111010010", -- 3537 FREE #<CONS 0 3538>
 "00000000000000000000110111010011", -- 3538 FREE #<CONS 0 3539>
 "00000000000000000000110111010100", -- 3539 FREE #<CONS 0 3540>
 "00000000000000000000110111010101", -- 3540 FREE #<CONS 0 3541>
 "00000000000000000000110111010110", -- 3541 FREE #<CONS 0 3542>
 "00000000000000000000110111010111", -- 3542 FREE #<CONS 0 3543>
 "00000000000000000000110111011000", -- 3543 FREE #<CONS 0 3544>
 "00000000000000000000110111011001", -- 3544 FREE #<CONS 0 3545>
 "00000000000000000000110111011010", -- 3545 FREE #<CONS 0 3546>
 "00000000000000000000110111011011", -- 3546 FREE #<CONS 0 3547>
 "00000000000000000000110111011100", -- 3547 FREE #<CONS 0 3548>
 "00000000000000000000110111011101", -- 3548 FREE #<CONS 0 3549>
 "00000000000000000000110111011110", -- 3549 FREE #<CONS 0 3550>
 "00000000000000000000110111011111", -- 3550 FREE #<CONS 0 3551>
 "00000000000000000000110111100000", -- 3551 FREE #<CONS 0 3552>
 "00000000000000000000110111100001", -- 3552 FREE #<CONS 0 3553>
 "00000000000000000000110111100010", -- 3553 FREE #<CONS 0 3554>
 "00000000000000000000110111100011", -- 3554 FREE #<CONS 0 3555>
 "00000000000000000000110111100100", -- 3555 FREE #<CONS 0 3556>
 "00000000000000000000110111100101", -- 3556 FREE #<CONS 0 3557>
 "00000000000000000000110111100110", -- 3557 FREE #<CONS 0 3558>
 "00000000000000000000110111100111", -- 3558 FREE #<CONS 0 3559>
 "00000000000000000000110111101000", -- 3559 FREE #<CONS 0 3560>
 "00000000000000000000110111101001", -- 3560 FREE #<CONS 0 3561>
 "00000000000000000000110111101010", -- 3561 FREE #<CONS 0 3562>
 "00000000000000000000110111101011", -- 3562 FREE #<CONS 0 3563>
 "00000000000000000000110111101100", -- 3563 FREE #<CONS 0 3564>
 "00000000000000000000110111101101", -- 3564 FREE #<CONS 0 3565>
 "00000000000000000000110111101110", -- 3565 FREE #<CONS 0 3566>
 "00000000000000000000110111101111", -- 3566 FREE #<CONS 0 3567>
 "00000000000000000000110111110000", -- 3567 FREE #<CONS 0 3568>
 "00000000000000000000110111110001", -- 3568 FREE #<CONS 0 3569>
 "00000000000000000000110111110010", -- 3569 FREE #<CONS 0 3570>
 "00000000000000000000110111110011", -- 3570 FREE #<CONS 0 3571>
 "00000000000000000000110111110100", -- 3571 FREE #<CONS 0 3572>
 "00000000000000000000110111110101", -- 3572 FREE #<CONS 0 3573>
 "00000000000000000000110111110110", -- 3573 FREE #<CONS 0 3574>
 "00000000000000000000110111110111", -- 3574 FREE #<CONS 0 3575>
 "00000000000000000000110111111000", -- 3575 FREE #<CONS 0 3576>
 "00000000000000000000110111111001", -- 3576 FREE #<CONS 0 3577>
 "00000000000000000000110111111010", -- 3577 FREE #<CONS 0 3578>
 "00000000000000000000110111111011", -- 3578 FREE #<CONS 0 3579>
 "00000000000000000000110111111100", -- 3579 FREE #<CONS 0 3580>
 "00000000000000000000110111111101", -- 3580 FREE #<CONS 0 3581>
 "00000000000000000000110111111110", -- 3581 FREE #<CONS 0 3582>
 "00000000000000000000110111111111", -- 3582 FREE #<CONS 0 3583>
 "00000000000000000000111000000000", -- 3583 FREE #<CONS 0 3584>
 "00000000000000000000111000000001", -- 3584 FREE #<CONS 0 3585>
 "00000000000000000000111000000010", -- 3585 FREE #<CONS 0 3586>
 "00000000000000000000111000000011", -- 3586 FREE #<CONS 0 3587>
 "00000000000000000000111000000100", -- 3587 FREE #<CONS 0 3588>
 "00000000000000000000111000000101", -- 3588 FREE #<CONS 0 3589>
 "00000000000000000000111000000110", -- 3589 FREE #<CONS 0 3590>
 "00000000000000000000111000000111", -- 3590 FREE #<CONS 0 3591>
 "00000000000000000000111000001000", -- 3591 FREE #<CONS 0 3592>
 "00000000000000000000111000001001", -- 3592 FREE #<CONS 0 3593>
 "00000000000000000000111000001010", -- 3593 FREE #<CONS 0 3594>
 "00000000000000000000111000001011", -- 3594 FREE #<CONS 0 3595>
 "00000000000000000000111000001100", -- 3595 FREE #<CONS 0 3596>
 "00000000000000000000111000001101", -- 3596 FREE #<CONS 0 3597>
 "00000000000000000000111000001110", -- 3597 FREE #<CONS 0 3598>
 "00000000000000000000111000001111", -- 3598 FREE #<CONS 0 3599>
 "00000000000000000000111000010000", -- 3599 FREE #<CONS 0 3600>
 "00000000000000000000111000010001", -- 3600 FREE #<CONS 0 3601>
 "00000000000000000000111000010010", -- 3601 FREE #<CONS 0 3602>
 "00000000000000000000111000010011", -- 3602 FREE #<CONS 0 3603>
 "00000000000000000000111000010100", -- 3603 FREE #<CONS 0 3604>
 "00000000000000000000111000010101", -- 3604 FREE #<CONS 0 3605>
 "00000000000000000000111000010110", -- 3605 FREE #<CONS 0 3606>
 "00000000000000000000111000010111", -- 3606 FREE #<CONS 0 3607>
 "00000000000000000000111000011000", -- 3607 FREE #<CONS 0 3608>
 "00000000000000000000111000011001", -- 3608 FREE #<CONS 0 3609>
 "00000000000000000000111000011010", -- 3609 FREE #<CONS 0 3610>
 "00000000000000000000111000011011", -- 3610 FREE #<CONS 0 3611>
 "00000000000000000000111000011100", -- 3611 FREE #<CONS 0 3612>
 "00000000000000000000111000011101", -- 3612 FREE #<CONS 0 3613>
 "00000000000000000000111000011110", -- 3613 FREE #<CONS 0 3614>
 "00000000000000000000111000011111", -- 3614 FREE #<CONS 0 3615>
 "00000000000000000000111000100000", -- 3615 FREE #<CONS 0 3616>
 "00000000000000000000111000100001", -- 3616 FREE #<CONS 0 3617>
 "00000000000000000000111000100010", -- 3617 FREE #<CONS 0 3618>
 "00000000000000000000111000100011", -- 3618 FREE #<CONS 0 3619>
 "00000000000000000000111000100100", -- 3619 FREE #<CONS 0 3620>
 "00000000000000000000111000100101", -- 3620 FREE #<CONS 0 3621>
 "00000000000000000000111000100110", -- 3621 FREE #<CONS 0 3622>
 "00000000000000000000111000100111", -- 3622 FREE #<CONS 0 3623>
 "00000000000000000000111000101000", -- 3623 FREE #<CONS 0 3624>
 "00000000000000000000111000101001", -- 3624 FREE #<CONS 0 3625>
 "00000000000000000000111000101010", -- 3625 FREE #<CONS 0 3626>
 "00000000000000000000111000101011", -- 3626 FREE #<CONS 0 3627>
 "00000000000000000000111000101100", -- 3627 FREE #<CONS 0 3628>
 "00000000000000000000111000101101", -- 3628 FREE #<CONS 0 3629>
 "00000000000000000000111000101110", -- 3629 FREE #<CONS 0 3630>
 "00000000000000000000111000101111", -- 3630 FREE #<CONS 0 3631>
 "00000000000000000000111000110000", -- 3631 FREE #<CONS 0 3632>
 "00000000000000000000111000110001", -- 3632 FREE #<CONS 0 3633>
 "00000000000000000000111000110010", -- 3633 FREE #<CONS 0 3634>
 "00000000000000000000111000110011", -- 3634 FREE #<CONS 0 3635>
 "00000000000000000000111000110100", -- 3635 FREE #<CONS 0 3636>
 "00000000000000000000111000110101", -- 3636 FREE #<CONS 0 3637>
 "00000000000000000000111000110110", -- 3637 FREE #<CONS 0 3638>
 "00000000000000000000111000110111", -- 3638 FREE #<CONS 0 3639>
 "00000000000000000000111000111000", -- 3639 FREE #<CONS 0 3640>
 "00000000000000000000111000111001", -- 3640 FREE #<CONS 0 3641>
 "00000000000000000000111000111010", -- 3641 FREE #<CONS 0 3642>
 "00000000000000000000111000111011", -- 3642 FREE #<CONS 0 3643>
 "00000000000000000000111000111100", -- 3643 FREE #<CONS 0 3644>
 "00000000000000000000111000111101", -- 3644 FREE #<CONS 0 3645>
 "00000000000000000000111000111110", -- 3645 FREE #<CONS 0 3646>
 "00000000000000000000111000111111", -- 3646 FREE #<CONS 0 3647>
 "00000000000000000000111001000000", -- 3647 FREE #<CONS 0 3648>
 "00000000000000000000111001000001", -- 3648 FREE #<CONS 0 3649>
 "00000000000000000000111001000010", -- 3649 FREE #<CONS 0 3650>
 "00000000000000000000111001000011", -- 3650 FREE #<CONS 0 3651>
 "00000000000000000000111001000100", -- 3651 FREE #<CONS 0 3652>
 "00000000000000000000111001000101", -- 3652 FREE #<CONS 0 3653>
 "00000000000000000000111001000110", -- 3653 FREE #<CONS 0 3654>
 "00000000000000000000111001000111", -- 3654 FREE #<CONS 0 3655>
 "00000000000000000000111001001000", -- 3655 FREE #<CONS 0 3656>
 "00000000000000000000111001001001", -- 3656 FREE #<CONS 0 3657>
 "00000000000000000000111001001010", -- 3657 FREE #<CONS 0 3658>
 "00000000000000000000111001001011", -- 3658 FREE #<CONS 0 3659>
 "00000000000000000000111001001100", -- 3659 FREE #<CONS 0 3660>
 "00000000000000000000111001001101", -- 3660 FREE #<CONS 0 3661>
 "00000000000000000000111001001110", -- 3661 FREE #<CONS 0 3662>
 "00000000000000000000111001001111", -- 3662 FREE #<CONS 0 3663>
 "00000000000000000000111001010000", -- 3663 FREE #<CONS 0 3664>
 "00000000000000000000111001010001", -- 3664 FREE #<CONS 0 3665>
 "00000000000000000000111001010010", -- 3665 FREE #<CONS 0 3666>
 "00000000000000000000111001010011", -- 3666 FREE #<CONS 0 3667>
 "00000000000000000000111001010100", -- 3667 FREE #<CONS 0 3668>
 "00000000000000000000111001010101", -- 3668 FREE #<CONS 0 3669>
 "00000000000000000000111001010110", -- 3669 FREE #<CONS 0 3670>
 "00000000000000000000111001010111", -- 3670 FREE #<CONS 0 3671>
 "00000000000000000000111001011000", -- 3671 FREE #<CONS 0 3672>
 "00000000000000000000111001011001", -- 3672 FREE #<CONS 0 3673>
 "00000000000000000000111001011010", -- 3673 FREE #<CONS 0 3674>
 "00000000000000000000111001011011", -- 3674 FREE #<CONS 0 3675>
 "00000000000000000000111001011100", -- 3675 FREE #<CONS 0 3676>
 "00000000000000000000111001011101", -- 3676 FREE #<CONS 0 3677>
 "00000000000000000000111001011110", -- 3677 FREE #<CONS 0 3678>
 "00000000000000000000111001011111", -- 3678 FREE #<CONS 0 3679>
 "00000000000000000000111001100000", -- 3679 FREE #<CONS 0 3680>
 "00000000000000000000111001100001", -- 3680 FREE #<CONS 0 3681>
 "00000000000000000000111001100010", -- 3681 FREE #<CONS 0 3682>
 "00000000000000000000111001100011", -- 3682 FREE #<CONS 0 3683>
 "00000000000000000000111001100100", -- 3683 FREE #<CONS 0 3684>
 "00000000000000000000111001100101", -- 3684 FREE #<CONS 0 3685>
 "00000000000000000000111001100110", -- 3685 FREE #<CONS 0 3686>
 "00000000000000000000111001100111", -- 3686 FREE #<CONS 0 3687>
 "00000000000000000000111001101000", -- 3687 FREE #<CONS 0 3688>
 "00000000000000000000111001101001", -- 3688 FREE #<CONS 0 3689>
 "00000000000000000000111001101010", -- 3689 FREE #<CONS 0 3690>
 "00000000000000000000111001101011", -- 3690 FREE #<CONS 0 3691>
 "00000000000000000000111001101100", -- 3691 FREE #<CONS 0 3692>
 "00000000000000000000111001101101", -- 3692 FREE #<CONS 0 3693>
 "00000000000000000000111001101110", -- 3693 FREE #<CONS 0 3694>
 "00000000000000000000111001101111", -- 3694 FREE #<CONS 0 3695>
 "00000000000000000000111001110000", -- 3695 FREE #<CONS 0 3696>
 "00000000000000000000111001110001", -- 3696 FREE #<CONS 0 3697>
 "00000000000000000000111001110010", -- 3697 FREE #<CONS 0 3698>
 "00000000000000000000111001110011", -- 3698 FREE #<CONS 0 3699>
 "00000000000000000000111001110100", -- 3699 FREE #<CONS 0 3700>
 "00000000000000000000111001110101", -- 3700 FREE #<CONS 0 3701>
 "00000000000000000000111001110110", -- 3701 FREE #<CONS 0 3702>
 "00000000000000000000111001110111", -- 3702 FREE #<CONS 0 3703>
 "00000000000000000000111001111000", -- 3703 FREE #<CONS 0 3704>
 "00000000000000000000111001111001", -- 3704 FREE #<CONS 0 3705>
 "00000000000000000000111001111010", -- 3705 FREE #<CONS 0 3706>
 "00000000000000000000111001111011", -- 3706 FREE #<CONS 0 3707>
 "00000000000000000000111001111100", -- 3707 FREE #<CONS 0 3708>
 "00000000000000000000111001111101", -- 3708 FREE #<CONS 0 3709>
 "00000000000000000000111001111110", -- 3709 FREE #<CONS 0 3710>
 "00000000000000000000111001111111", -- 3710 FREE #<CONS 0 3711>
 "00000000000000000000111010000000", -- 3711 FREE #<CONS 0 3712>
 "00000000000000000000111010000001", -- 3712 FREE #<CONS 0 3713>
 "00000000000000000000111010000010", -- 3713 FREE #<CONS 0 3714>
 "00000000000000000000111010000011", -- 3714 FREE #<CONS 0 3715>
 "00000000000000000000111010000100", -- 3715 FREE #<CONS 0 3716>
 "00000000000000000000111010000101", -- 3716 FREE #<CONS 0 3717>
 "00000000000000000000111010000110", -- 3717 FREE #<CONS 0 3718>
 "00000000000000000000111010000111", -- 3718 FREE #<CONS 0 3719>
 "00000000000000000000111010001000", -- 3719 FREE #<CONS 0 3720>
 "00000000000000000000111010001001", -- 3720 FREE #<CONS 0 3721>
 "00000000000000000000111010001010", -- 3721 FREE #<CONS 0 3722>
 "00000000000000000000111010001011", -- 3722 FREE #<CONS 0 3723>
 "00000000000000000000111010001100", -- 3723 FREE #<CONS 0 3724>
 "00000000000000000000111010001101", -- 3724 FREE #<CONS 0 3725>
 "00000000000000000000111010001110", -- 3725 FREE #<CONS 0 3726>
 "00000000000000000000111010001111", -- 3726 FREE #<CONS 0 3727>
 "00000000000000000000111010010000", -- 3727 FREE #<CONS 0 3728>
 "00000000000000000000111010010001", -- 3728 FREE #<CONS 0 3729>
 "00000000000000000000111010010010", -- 3729 FREE #<CONS 0 3730>
 "00000000000000000000111010010011", -- 3730 FREE #<CONS 0 3731>
 "00000000000000000000111010010100", -- 3731 FREE #<CONS 0 3732>
 "00000000000000000000111010010101", -- 3732 FREE #<CONS 0 3733>
 "00000000000000000000111010010110", -- 3733 FREE #<CONS 0 3734>
 "00000000000000000000111010010111", -- 3734 FREE #<CONS 0 3735>
 "00000000000000000000111010011000", -- 3735 FREE #<CONS 0 3736>
 "00000000000000000000111010011001", -- 3736 FREE #<CONS 0 3737>
 "00000000000000000000111010011010", -- 3737 FREE #<CONS 0 3738>
 "00000000000000000000111010011011", -- 3738 FREE #<CONS 0 3739>
 "00000000000000000000111010011100", -- 3739 FREE #<CONS 0 3740>
 "00000000000000000000111010011101", -- 3740 FREE #<CONS 0 3741>
 "00000000000000000000111010011110", -- 3741 FREE #<CONS 0 3742>
 "00000000000000000000111010011111", -- 3742 FREE #<CONS 0 3743>
 "00000000000000000000111010100000", -- 3743 FREE #<CONS 0 3744>
 "00000000000000000000111010100001", -- 3744 FREE #<CONS 0 3745>
 "00000000000000000000111010100010", -- 3745 FREE #<CONS 0 3746>
 "00000000000000000000111010100011", -- 3746 FREE #<CONS 0 3747>
 "00000000000000000000111010100100", -- 3747 FREE #<CONS 0 3748>
 "00000000000000000000111010100101", -- 3748 FREE #<CONS 0 3749>
 "00000000000000000000111010100110", -- 3749 FREE #<CONS 0 3750>
 "00000000000000000000111010100111", -- 3750 FREE #<CONS 0 3751>
 "00000000000000000000111010101000", -- 3751 FREE #<CONS 0 3752>
 "00000000000000000000111010101001", -- 3752 FREE #<CONS 0 3753>
 "00000000000000000000111010101010", -- 3753 FREE #<CONS 0 3754>
 "00000000000000000000111010101011", -- 3754 FREE #<CONS 0 3755>
 "00000000000000000000111010101100", -- 3755 FREE #<CONS 0 3756>
 "00000000000000000000111010101101", -- 3756 FREE #<CONS 0 3757>
 "00000000000000000000111010101110", -- 3757 FREE #<CONS 0 3758>
 "00000000000000000000111010101111", -- 3758 FREE #<CONS 0 3759>
 "00000000000000000000111010110000", -- 3759 FREE #<CONS 0 3760>
 "00000000000000000000111010110001", -- 3760 FREE #<CONS 0 3761>
 "00000000000000000000111010110010", -- 3761 FREE #<CONS 0 3762>
 "00000000000000000000111010110011", -- 3762 FREE #<CONS 0 3763>
 "00000000000000000000111010110100", -- 3763 FREE #<CONS 0 3764>
 "00000000000000000000111010110101", -- 3764 FREE #<CONS 0 3765>
 "00000000000000000000111010110110", -- 3765 FREE #<CONS 0 3766>
 "00000000000000000000111010110111", -- 3766 FREE #<CONS 0 3767>
 "00000000000000000000111010111000", -- 3767 FREE #<CONS 0 3768>
 "00000000000000000000111010111001", -- 3768 FREE #<CONS 0 3769>
 "00000000000000000000111010111010", -- 3769 FREE #<CONS 0 3770>
 "00000000000000000000111010111011", -- 3770 FREE #<CONS 0 3771>
 "00000000000000000000111010111100", -- 3771 FREE #<CONS 0 3772>
 "00000000000000000000111010111101", -- 3772 FREE #<CONS 0 3773>
 "00000000000000000000111010111110", -- 3773 FREE #<CONS 0 3774>
 "00000000000000000000111010111111", -- 3774 FREE #<CONS 0 3775>
 "00000000000000000000111011000000", -- 3775 FREE #<CONS 0 3776>
 "00000000000000000000111011000001", -- 3776 FREE #<CONS 0 3777>
 "00000000000000000000111011000010", -- 3777 FREE #<CONS 0 3778>
 "00000000000000000000111011000011", -- 3778 FREE #<CONS 0 3779>
 "00000000000000000000111011000100", -- 3779 FREE #<CONS 0 3780>
 "00000000000000000000111011000101", -- 3780 FREE #<CONS 0 3781>
 "00000000000000000000111011000110", -- 3781 FREE #<CONS 0 3782>
 "00000000000000000000111011000111", -- 3782 FREE #<CONS 0 3783>
 "00000000000000000000111011001000", -- 3783 FREE #<CONS 0 3784>
 "00000000000000000000111011001001", -- 3784 FREE #<CONS 0 3785>
 "00000000000000000000111011001010", -- 3785 FREE #<CONS 0 3786>
 "00000000000000000000111011001011", -- 3786 FREE #<CONS 0 3787>
 "00000000000000000000111011001100", -- 3787 FREE #<CONS 0 3788>
 "00000000000000000000111011001101", -- 3788 FREE #<CONS 0 3789>
 "00000000000000000000111011001110", -- 3789 FREE #<CONS 0 3790>
 "00000000000000000000111011001111", -- 3790 FREE #<CONS 0 3791>
 "00000000000000000000111011010000", -- 3791 FREE #<CONS 0 3792>
 "00000000000000000000111011010001", -- 3792 FREE #<CONS 0 3793>
 "00000000000000000000111011010010", -- 3793 FREE #<CONS 0 3794>
 "00000000000000000000111011010011", -- 3794 FREE #<CONS 0 3795>
 "00000000000000000000111011010100", -- 3795 FREE #<CONS 0 3796>
 "00000000000000000000111011010101", -- 3796 FREE #<CONS 0 3797>
 "00000000000000000000111011010110", -- 3797 FREE #<CONS 0 3798>
 "00000000000000000000111011010111", -- 3798 FREE #<CONS 0 3799>
 "00000000000000000000111011011000", -- 3799 FREE #<CONS 0 3800>
 "00000000000000000000111011011001", -- 3800 FREE #<CONS 0 3801>
 "00000000000000000000111011011010", -- 3801 FREE #<CONS 0 3802>
 "00000000000000000000111011011011", -- 3802 FREE #<CONS 0 3803>
 "00000000000000000000111011011100", -- 3803 FREE #<CONS 0 3804>
 "00000000000000000000111011011101", -- 3804 FREE #<CONS 0 3805>
 "00000000000000000000111011011110", -- 3805 FREE #<CONS 0 3806>
 "00000000000000000000111011011111", -- 3806 FREE #<CONS 0 3807>
 "00000000000000000000111011100000", -- 3807 FREE #<CONS 0 3808>
 "00000000000000000000111011100001", -- 3808 FREE #<CONS 0 3809>
 "00000000000000000000111011100010", -- 3809 FREE #<CONS 0 3810>
 "00000000000000000000111011100011", -- 3810 FREE #<CONS 0 3811>
 "00000000000000000000111011100100", -- 3811 FREE #<CONS 0 3812>
 "00000000000000000000111011100101", -- 3812 FREE #<CONS 0 3813>
 "00000000000000000000111011100110", -- 3813 FREE #<CONS 0 3814>
 "00000000000000000000111011100111", -- 3814 FREE #<CONS 0 3815>
 "00000000000000000000111011101000", -- 3815 FREE #<CONS 0 3816>
 "00000000000000000000111011101001", -- 3816 FREE #<CONS 0 3817>
 "00000000000000000000111011101010", -- 3817 FREE #<CONS 0 3818>
 "00000000000000000000111011101011", -- 3818 FREE #<CONS 0 3819>
 "00000000000000000000111011101100", -- 3819 FREE #<CONS 0 3820>
 "00000000000000000000111011101101", -- 3820 FREE #<CONS 0 3821>
 "00000000000000000000111011101110", -- 3821 FREE #<CONS 0 3822>
 "00000000000000000000111011101111", -- 3822 FREE #<CONS 0 3823>
 "00000000000000000000111011110000", -- 3823 FREE #<CONS 0 3824>
 "00000000000000000000111011110001", -- 3824 FREE #<CONS 0 3825>
 "00000000000000000000111011110010", -- 3825 FREE #<CONS 0 3826>
 "00000000000000000000111011110011", -- 3826 FREE #<CONS 0 3827>
 "00000000000000000000111011110100", -- 3827 FREE #<CONS 0 3828>
 "00000000000000000000111011110101", -- 3828 FREE #<CONS 0 3829>
 "00000000000000000000111011110110", -- 3829 FREE #<CONS 0 3830>
 "00000000000000000000111011110111", -- 3830 FREE #<CONS 0 3831>
 "00000000000000000000111011111000", -- 3831 FREE #<CONS 0 3832>
 "00000000000000000000111011111001", -- 3832 FREE #<CONS 0 3833>
 "00000000000000000000111011111010", -- 3833 FREE #<CONS 0 3834>
 "00000000000000000000111011111011", -- 3834 FREE #<CONS 0 3835>
 "00000000000000000000111011111100", -- 3835 FREE #<CONS 0 3836>
 "00000000000000000000111011111101", -- 3836 FREE #<CONS 0 3837>
 "00000000000000000000111011111110", -- 3837 FREE #<CONS 0 3838>
 "00000000000000000000111011111111", -- 3838 FREE #<CONS 0 3839>
 "00000000000000000000111100000000", -- 3839 FREE #<CONS 0 3840>
 "00000000000000000000111100000001", -- 3840 FREE #<CONS 0 3841>
 "00000000000000000000111100000010", -- 3841 FREE #<CONS 0 3842>
 "00000000000000000000111100000011", -- 3842 FREE #<CONS 0 3843>
 "00000000000000000000111100000100", -- 3843 FREE #<CONS 0 3844>
 "00000000000000000000111100000101", -- 3844 FREE #<CONS 0 3845>
 "00000000000000000000111100000110", -- 3845 FREE #<CONS 0 3846>
 "00000000000000000000111100000111", -- 3846 FREE #<CONS 0 3847>
 "00000000000000000000111100001000", -- 3847 FREE #<CONS 0 3848>
 "00000000000000000000111100001001", -- 3848 FREE #<CONS 0 3849>
 "00000000000000000000111100001010", -- 3849 FREE #<CONS 0 3850>
 "00000000000000000000111100001011", -- 3850 FREE #<CONS 0 3851>
 "00000000000000000000111100001100", -- 3851 FREE #<CONS 0 3852>
 "00000000000000000000111100001101", -- 3852 FREE #<CONS 0 3853>
 "00000000000000000000111100001110", -- 3853 FREE #<CONS 0 3854>
 "00000000000000000000111100001111", -- 3854 FREE #<CONS 0 3855>
 "00000000000000000000111100010000", -- 3855 FREE #<CONS 0 3856>
 "00000000000000000000111100010001", -- 3856 FREE #<CONS 0 3857>
 "00000000000000000000111100010010", -- 3857 FREE #<CONS 0 3858>
 "00000000000000000000111100010011", -- 3858 FREE #<CONS 0 3859>
 "00000000000000000000111100010100", -- 3859 FREE #<CONS 0 3860>
 "00000000000000000000111100010101", -- 3860 FREE #<CONS 0 3861>
 "00000000000000000000111100010110", -- 3861 FREE #<CONS 0 3862>
 "00000000000000000000111100010111", -- 3862 FREE #<CONS 0 3863>
 "00000000000000000000111100011000", -- 3863 FREE #<CONS 0 3864>
 "00000000000000000000111100011001", -- 3864 FREE #<CONS 0 3865>
 "00000000000000000000111100011010", -- 3865 FREE #<CONS 0 3866>
 "00000000000000000000111100011011", -- 3866 FREE #<CONS 0 3867>
 "00000000000000000000111100011100", -- 3867 FREE #<CONS 0 3868>
 "00000000000000000000111100011101", -- 3868 FREE #<CONS 0 3869>
 "00000000000000000000111100011110", -- 3869 FREE #<CONS 0 3870>
 "00000000000000000000111100011111", -- 3870 FREE #<CONS 0 3871>
 "00000000000000000000111100100000", -- 3871 FREE #<CONS 0 3872>
 "00000000000000000000111100100001", -- 3872 FREE #<CONS 0 3873>
 "00000000000000000000111100100010", -- 3873 FREE #<CONS 0 3874>
 "00000000000000000000111100100011", -- 3874 FREE #<CONS 0 3875>
 "00000000000000000000111100100100", -- 3875 FREE #<CONS 0 3876>
 "00000000000000000000111100100101", -- 3876 FREE #<CONS 0 3877>
 "00000000000000000000111100100110", -- 3877 FREE #<CONS 0 3878>
 "00000000000000000000111100100111", -- 3878 FREE #<CONS 0 3879>
 "00000000000000000000111100101000", -- 3879 FREE #<CONS 0 3880>
 "00000000000000000000111100101001", -- 3880 FREE #<CONS 0 3881>
 "00000000000000000000111100101010", -- 3881 FREE #<CONS 0 3882>
 "00000000000000000000111100101011", -- 3882 FREE #<CONS 0 3883>
 "00000000000000000000111100101100", -- 3883 FREE #<CONS 0 3884>
 "00000000000000000000111100101101", -- 3884 FREE #<CONS 0 3885>
 "00000000000000000000111100101110", -- 3885 FREE #<CONS 0 3886>
 "00000000000000000000111100101111", -- 3886 FREE #<CONS 0 3887>
 "00000000000000000000111100110000", -- 3887 FREE #<CONS 0 3888>
 "00000000000000000000111100110001", -- 3888 FREE #<CONS 0 3889>
 "00000000000000000000111100110010", -- 3889 FREE #<CONS 0 3890>
 "00000000000000000000111100110011", -- 3890 FREE #<CONS 0 3891>
 "00000000000000000000111100110100", -- 3891 FREE #<CONS 0 3892>
 "00000000000000000000111100110101", -- 3892 FREE #<CONS 0 3893>
 "00000000000000000000111100110110", -- 3893 FREE #<CONS 0 3894>
 "00000000000000000000111100110111", -- 3894 FREE #<CONS 0 3895>
 "00000000000000000000111100111000", -- 3895 FREE #<CONS 0 3896>
 "00000000000000000000111100111001", -- 3896 FREE #<CONS 0 3897>
 "00000000000000000000111100111010", -- 3897 FREE #<CONS 0 3898>
 "00000000000000000000111100111011", -- 3898 FREE #<CONS 0 3899>
 "00000000000000000000111100111100", -- 3899 FREE #<CONS 0 3900>
 "00000000000000000000111100111101", -- 3900 FREE #<CONS 0 3901>
 "00000000000000000000111100111110", -- 3901 FREE #<CONS 0 3902>
 "00000000000000000000111100111111", -- 3902 FREE #<CONS 0 3903>
 "00000000000000000000111101000000", -- 3903 FREE #<CONS 0 3904>
 "00000000000000000000111101000001", -- 3904 FREE #<CONS 0 3905>
 "00000000000000000000111101000010", -- 3905 FREE #<CONS 0 3906>
 "00000000000000000000111101000011", -- 3906 FREE #<CONS 0 3907>
 "00000000000000000000111101000100", -- 3907 FREE #<CONS 0 3908>
 "00000000000000000000111101000101", -- 3908 FREE #<CONS 0 3909>
 "00000000000000000000111101000110", -- 3909 FREE #<CONS 0 3910>
 "00000000000000000000111101000111", -- 3910 FREE #<CONS 0 3911>
 "00000000000000000000111101001000", -- 3911 FREE #<CONS 0 3912>
 "00000000000000000000111101001001", -- 3912 FREE #<CONS 0 3913>
 "00000000000000000000111101001010", -- 3913 FREE #<CONS 0 3914>
 "00000000000000000000111101001011", -- 3914 FREE #<CONS 0 3915>
 "00000000000000000000111101001100", -- 3915 FREE #<CONS 0 3916>
 "00000000000000000000111101001101", -- 3916 FREE #<CONS 0 3917>
 "00000000000000000000111101001110", -- 3917 FREE #<CONS 0 3918>
 "00000000000000000000111101001111", -- 3918 FREE #<CONS 0 3919>
 "00000000000000000000111101010000", -- 3919 FREE #<CONS 0 3920>
 "00000000000000000000111101010001", -- 3920 FREE #<CONS 0 3921>
 "00000000000000000000111101010010", -- 3921 FREE #<CONS 0 3922>
 "00000000000000000000111101010011", -- 3922 FREE #<CONS 0 3923>
 "00000000000000000000111101010100", -- 3923 FREE #<CONS 0 3924>
 "00000000000000000000111101010101", -- 3924 FREE #<CONS 0 3925>
 "00000000000000000000111101010110", -- 3925 FREE #<CONS 0 3926>
 "00000000000000000000111101010111", -- 3926 FREE #<CONS 0 3927>
 "00000000000000000000111101011000", -- 3927 FREE #<CONS 0 3928>
 "00000000000000000000111101011001", -- 3928 FREE #<CONS 0 3929>
 "00000000000000000000111101011010", -- 3929 FREE #<CONS 0 3930>
 "00000000000000000000111101011011", -- 3930 FREE #<CONS 0 3931>
 "00000000000000000000111101011100", -- 3931 FREE #<CONS 0 3932>
 "00000000000000000000111101011101", -- 3932 FREE #<CONS 0 3933>
 "00000000000000000000111101011110", -- 3933 FREE #<CONS 0 3934>
 "00000000000000000000111101011111", -- 3934 FREE #<CONS 0 3935>
 "00000000000000000000111101100000", -- 3935 FREE #<CONS 0 3936>
 "00000000000000000000111101100001", -- 3936 FREE #<CONS 0 3937>
 "00000000000000000000111101100010", -- 3937 FREE #<CONS 0 3938>
 "00000000000000000000111101100011", -- 3938 FREE #<CONS 0 3939>
 "00000000000000000000111101100100", -- 3939 FREE #<CONS 0 3940>
 "00000000000000000000111101100101", -- 3940 FREE #<CONS 0 3941>
 "00000000000000000000111101100110", -- 3941 FREE #<CONS 0 3942>
 "00000000000000000000111101100111", -- 3942 FREE #<CONS 0 3943>
 "00000000000000000000111101101000", -- 3943 FREE #<CONS 0 3944>
 "00000000000000000000111101101001", -- 3944 FREE #<CONS 0 3945>
 "00000000000000000000111101101010", -- 3945 FREE #<CONS 0 3946>
 "00000000000000000000111101101011", -- 3946 FREE #<CONS 0 3947>
 "00000000000000000000111101101100", -- 3947 FREE #<CONS 0 3948>
 "00000000000000000000111101101101", -- 3948 FREE #<CONS 0 3949>
 "00000000000000000000111101101110", -- 3949 FREE #<CONS 0 3950>
 "00000000000000000000111101101111", -- 3950 FREE #<CONS 0 3951>
 "00000000000000000000111101110000", -- 3951 FREE #<CONS 0 3952>
 "00000000000000000000111101110001", -- 3952 FREE #<CONS 0 3953>
 "00000000000000000000111101110010", -- 3953 FREE #<CONS 0 3954>
 "00000000000000000000111101110011", -- 3954 FREE #<CONS 0 3955>
 "00000000000000000000111101110100", -- 3955 FREE #<CONS 0 3956>
 "00000000000000000000111101110101", -- 3956 FREE #<CONS 0 3957>
 "00000000000000000000111101110110", -- 3957 FREE #<CONS 0 3958>
 "00000000000000000000111101110111", -- 3958 FREE #<CONS 0 3959>
 "00000000000000000000111101111000", -- 3959 FREE #<CONS 0 3960>
 "00000000000000000000111101111001", -- 3960 FREE #<CONS 0 3961>
 "00000000000000000000111101111010", -- 3961 FREE #<CONS 0 3962>
 "00000000000000000000111101111011", -- 3962 FREE #<CONS 0 3963>
 "00000000000000000000111101111100", -- 3963 FREE #<CONS 0 3964>
 "00000000000000000000111101111101", -- 3964 FREE #<CONS 0 3965>
 "00000000000000000000111101111110", -- 3965 FREE #<CONS 0 3966>
 "00000000000000000000111101111111", -- 3966 FREE #<CONS 0 3967>
 "00000000000000000000111110000000", -- 3967 FREE #<CONS 0 3968>
 "00000000000000000000111110000001", -- 3968 FREE #<CONS 0 3969>
 "00000000000000000000111110000010", -- 3969 FREE #<CONS 0 3970>
 "00000000000000000000111110000011", -- 3970 FREE #<CONS 0 3971>
 "00000000000000000000111110000100", -- 3971 FREE #<CONS 0 3972>
 "00000000000000000000111110000101", -- 3972 FREE #<CONS 0 3973>
 "00000000000000000000111110000110", -- 3973 FREE #<CONS 0 3974>
 "00000000000000000000111110000111", -- 3974 FREE #<CONS 0 3975>
 "00000000000000000000111110001000", -- 3975 FREE #<CONS 0 3976>
 "00000000000000000000111110001001", -- 3976 FREE #<CONS 0 3977>
 "00000000000000000000111110001010", -- 3977 FREE #<CONS 0 3978>
 "00000000000000000000111110001011", -- 3978 FREE #<CONS 0 3979>
 "00000000000000000000111110001100", -- 3979 FREE #<CONS 0 3980>
 "00000000000000000000111110001101", -- 3980 FREE #<CONS 0 3981>
 "00000000000000000000111110001110", -- 3981 FREE #<CONS 0 3982>
 "00000000000000000000111110001111", -- 3982 FREE #<CONS 0 3983>
 "00000000000000000000111110010000", -- 3983 FREE #<CONS 0 3984>
 "00000000000000000000111110010001", -- 3984 FREE #<CONS 0 3985>
 "00000000000000000000111110010010", -- 3985 FREE #<CONS 0 3986>
 "00000000000000000000111110010011", -- 3986 FREE #<CONS 0 3987>
 "00000000000000000000111110010100", -- 3987 FREE #<CONS 0 3988>
 "00000000000000000000111110010101", -- 3988 FREE #<CONS 0 3989>
 "00000000000000000000111110010110", -- 3989 FREE #<CONS 0 3990>
 "00000000000000000000111110010111", -- 3990 FREE #<CONS 0 3991>
 "00000000000000000000111110011000", -- 3991 FREE #<CONS 0 3992>
 "00000000000000000000111110011001", -- 3992 FREE #<CONS 0 3993>
 "00000000000000000000111110011010", -- 3993 FREE #<CONS 0 3994>
 "00000000000000000000111110011011", -- 3994 FREE #<CONS 0 3995>
 "00000000000000000000111110011100", -- 3995 FREE #<CONS 0 3996>
 "00000000000000000000111110011101", -- 3996 FREE #<CONS 0 3997>
 "00000000000000000000111110011110", -- 3997 FREE #<CONS 0 3998>
 "00000000000000000000111110011111", -- 3998 FREE #<CONS 0 3999>
 "00000000000000000000111110100000", -- 3999 FREE #<CONS 0 4000>
 "00000000000000000000111110100001", -- 4000 FREE #<CONS 0 4001>
 "00000000000000000000111110100010", -- 4001 FREE #<CONS 0 4002>
 "00000000000000000000111110100011", -- 4002 FREE #<CONS 0 4003>
 "00000000000000000000111110100100", -- 4003 FREE #<CONS 0 4004>
 "00000000000000000000111110100101", -- 4004 FREE #<CONS 0 4005>
 "00000000000000000000111110100110", -- 4005 FREE #<CONS 0 4006>
 "00000000000000000000111110100111", -- 4006 FREE #<CONS 0 4007>
 "00000000000000000000111110101000", -- 4007 FREE #<CONS 0 4008>
 "00000000000000000000111110101001", -- 4008 FREE #<CONS 0 4009>
 "00000000000000000000111110101010", -- 4009 FREE #<CONS 0 4010>
 "00000000000000000000111110101011", -- 4010 FREE #<CONS 0 4011>
 "00000000000000000000111110101100", -- 4011 FREE #<CONS 0 4012>
 "00000000000000000000111110101101", -- 4012 FREE #<CONS 0 4013>
 "00000000000000000000111110101110", -- 4013 FREE #<CONS 0 4014>
 "00000000000000000000111110101111", -- 4014 FREE #<CONS 0 4015>
 "00000000000000000000111110110000", -- 4015 FREE #<CONS 0 4016>
 "00000000000000000000111110110001", -- 4016 FREE #<CONS 0 4017>
 "00000000000000000000111110110010", -- 4017 FREE #<CONS 0 4018>
 "00000000000000000000111110110011", -- 4018 FREE #<CONS 0 4019>
 "00000000000000000000111110110100", -- 4019 FREE #<CONS 0 4020>
 "00000000000000000000111110110101", -- 4020 FREE #<CONS 0 4021>
 "00000000000000000000111110110110", -- 4021 FREE #<CONS 0 4022>
 "00000000000000000000111110110111", -- 4022 FREE #<CONS 0 4023>
 "00000000000000000000111110111000", -- 4023 FREE #<CONS 0 4024>
 "00000000000000000000111110111001", -- 4024 FREE #<CONS 0 4025>
 "00000000000000000000111110111010", -- 4025 FREE #<CONS 0 4026>
 "00000000000000000000111110111011", -- 4026 FREE #<CONS 0 4027>
 "00000000000000000000111110111100", -- 4027 FREE #<CONS 0 4028>
 "00000000000000000000111110111101", -- 4028 FREE #<CONS 0 4029>
 "00000000000000000000111110111110", -- 4029 FREE #<CONS 0 4030>
 "00000000000000000000111110111111", -- 4030 FREE #<CONS 0 4031>
 "00000000000000000000111111000000", -- 4031 FREE #<CONS 0 4032>
 "00000000000000000000111111000001", -- 4032 FREE #<CONS 0 4033>
 "00000000000000000000111111000010", -- 4033 FREE #<CONS 0 4034>
 "00000000000000000000111111000011", -- 4034 FREE #<CONS 0 4035>
 "00000000000000000000111111000100", -- 4035 FREE #<CONS 0 4036>
 "00000000000000000000111111000101", -- 4036 FREE #<CONS 0 4037>
 "00000000000000000000111111000110", -- 4037 FREE #<CONS 0 4038>
 "00000000000000000000111111000111", -- 4038 FREE #<CONS 0 4039>
 "00000000000000000000111111001000", -- 4039 FREE #<CONS 0 4040>
 "00000000000000000000111111001001", -- 4040 FREE #<CONS 0 4041>
 "00000000000000000000111111001010", -- 4041 FREE #<CONS 0 4042>
 "00000000000000000000111111001011", -- 4042 FREE #<CONS 0 4043>
 "00000000000000000000111111001100", -- 4043 FREE #<CONS 0 4044>
 "00000000000000000000111111001101", -- 4044 FREE #<CONS 0 4045>
 "00000000000000000000111111001110", -- 4045 FREE #<CONS 0 4046>
 "00000000000000000000111111001111", -- 4046 FREE #<CONS 0 4047>
 "00000000000000000000111111010000", -- 4047 FREE #<CONS 0 4048>
 "00000000000000000000111111010001", -- 4048 FREE #<CONS 0 4049>
 "00000000000000000000111111010010", -- 4049 FREE #<CONS 0 4050>
 "00000000000000000000111111010011", -- 4050 FREE #<CONS 0 4051>
 "00000000000000000000111111010100", -- 4051 FREE #<CONS 0 4052>
 "00000000000000000000111111010101", -- 4052 FREE #<CONS 0 4053>
 "00000000000000000000111111010110", -- 4053 FREE #<CONS 0 4054>
 "00000000000000000000111111010111", -- 4054 FREE #<CONS 0 4055>
 "00000000000000000000111111011000", -- 4055 FREE #<CONS 0 4056>
 "00000000000000000000111111011001", -- 4056 FREE #<CONS 0 4057>
 "00000000000000000000111111011010", -- 4057 FREE #<CONS 0 4058>
 "00000000000000000000111111011011", -- 4058 FREE #<CONS 0 4059>
 "00000000000000000000111111011100", -- 4059 FREE #<CONS 0 4060>
 "00000000000000000000111111011101", -- 4060 FREE #<CONS 0 4061>
 "00000000000000000000111111011110", -- 4061 FREE #<CONS 0 4062>
 "00000000000000000000111111011111", -- 4062 FREE #<CONS 0 4063>
 "00000000000000000000111111100000", -- 4063 FREE #<CONS 0 4064>
 "00000000000000000000111111100001", -- 4064 FREE #<CONS 0 4065>
 "00000000000000000000111111100010", -- 4065 FREE #<CONS 0 4066>
 "00000000000000000000111111100011", -- 4066 FREE #<CONS 0 4067>
 "00000000000000000000111111100100", -- 4067 FREE #<CONS 0 4068>
 "00000000000000000000111111100101", -- 4068 FREE #<CONS 0 4069>
 "00000000000000000000111111100110", -- 4069 FREE #<CONS 0 4070>
 "00000000000000000000111111100111", -- 4070 FREE #<CONS 0 4071>
 "00000000000000000000111111101000", -- 4071 FREE #<CONS 0 4072>
 "00000000000000000000111111101001", -- 4072 FREE #<CONS 0 4073>
 "00000000000000000000111111101010", -- 4073 FREE #<CONS 0 4074>
 "00000000000000000000111111101011", -- 4074 FREE #<CONS 0 4075>
 "00000000000000000000111111101100", -- 4075 FREE #<CONS 0 4076>
 "00000000000000000000111111101101", -- 4076 FREE #<CONS 0 4077>
 "00000000000000000000111111101110", -- 4077 FREE #<CONS 0 4078>
 "00000000000000000000111111101111", -- 4078 FREE #<CONS 0 4079>
 "00000000000000000000111111110000", -- 4079 FREE #<CONS 0 4080>
 "00000000000000000000111111110001", -- 4080 FREE #<CONS 0 4081>
 "00000000000000000000111111110010", -- 4081 FREE #<CONS 0 4082>
 "00000000000000000000111111110011", -- 4082 FREE #<CONS 0 4083>
 "00000000000000000000111111110100", -- 4083 FREE #<CONS 0 4084>
 "00000000000000000000111111110101", -- 4084 FREE #<CONS 0 4085>
 "00000000000000000000111111110110", -- 4085 FREE #<CONS 0 4086>
 "00000000000000000000111111110111", -- 4086 FREE #<CONS 0 4087>
 "00000000000000000000111111111000", -- 4087 FREE #<CONS 0 4088>
 "00000000000000000000111111111001", -- 4088 FREE #<CONS 0 4089>
 "00000000000000000000111111111010", -- 4089 FREE #<CONS 0 4090>
 "00000000000000000000111111111011", -- 4090 FREE #<CONS 0 4091>
 "00000000000000000000111111111100", -- 4091 FREE #<CONS 0 4092>
 "00000000000000000000111111111101", -- 4092 FREE #<CONS 0 4093>
 "00000000000000000000111111111110", -- 4093 FREE #<CONS 0 4094>
 "00000000000000000000111111111111", -- 4094 FREE #<CONS 0 4095>
 "00000000000000000001000000000000", -- 4095 FREE #<CONS 0 4096>
 "00000000000000000001000000000001", -- 4096 FREE #<CONS 0 4097>
 "00000000000000000001000000000010", -- 4097 FREE #<CONS 0 4098>
 "00000000000000000001000000000011", -- 4098 FREE #<CONS 0 4099>
 "00000000000000000001000000000100", -- 4099 FREE #<CONS 0 4100>
 "00000000000000000001000000000101", -- 4100 FREE #<CONS 0 4101>
 "00000000000000000001000000000110", -- 4101 FREE #<CONS 0 4102>
 "00000000000000000001000000000111", -- 4102 FREE #<CONS 0 4103>
 "00000000000000000001000000001000", -- 4103 FREE #<CONS 0 4104>
 "00000000000000000001000000001001", -- 4104 FREE #<CONS 0 4105>
 "00000000000000000001000000001010", -- 4105 FREE #<CONS 0 4106>
 "00000000000000000001000000001011", -- 4106 FREE #<CONS 0 4107>
 "00000000000000000001000000001100", -- 4107 FREE #<CONS 0 4108>
 "00000000000000000001000000001101", -- 4108 FREE #<CONS 0 4109>
 "00000000000000000001000000001110", -- 4109 FREE #<CONS 0 4110>
 "00000000000000000001000000001111", -- 4110 FREE #<CONS 0 4111>
 "00000000000000000001000000010000", -- 4111 FREE #<CONS 0 4112>
 "00000000000000000001000000010001", -- 4112 FREE #<CONS 0 4113>
 "00000000000000000001000000010010", -- 4113 FREE #<CONS 0 4114>
 "00000000000000000001000000010011", -- 4114 FREE #<CONS 0 4115>
 "00000000000000000001000000010100", -- 4115 FREE #<CONS 0 4116>
 "00000000000000000001000000010101", -- 4116 FREE #<CONS 0 4117>
 "00000000000000000001000000010110", -- 4117 FREE #<CONS 0 4118>
 "00000000000000000001000000010111", -- 4118 FREE #<CONS 0 4119>
 "00000000000000000001000000011000", -- 4119 FREE #<CONS 0 4120>
 "00000000000000000001000000011001", -- 4120 FREE #<CONS 0 4121>
 "00000000000000000001000000011010", -- 4121 FREE #<CONS 0 4122>
 "00000000000000000001000000011011", -- 4122 FREE #<CONS 0 4123>
 "00000000000000000001000000011100", -- 4123 FREE #<CONS 0 4124>
 "00000000000000000001000000011101", -- 4124 FREE #<CONS 0 4125>
 "00000000000000000001000000011110", -- 4125 FREE #<CONS 0 4126>
 "00000000000000000001000000011111", -- 4126 FREE #<CONS 0 4127>
 "00000000000000000001000000100000", -- 4127 FREE #<CONS 0 4128>
 "00000000000000000001000000100001", -- 4128 FREE #<CONS 0 4129>
 "00000000000000000001000000100010", -- 4129 FREE #<CONS 0 4130>
 "00000000000000000001000000100011", -- 4130 FREE #<CONS 0 4131>
 "00000000000000000001000000100100", -- 4131 FREE #<CONS 0 4132>
 "00000000000000000001000000100101", -- 4132 FREE #<CONS 0 4133>
 "00000000000000000001000000100110", -- 4133 FREE #<CONS 0 4134>
 "00000000000000000001000000100111", -- 4134 FREE #<CONS 0 4135>
 "00000000000000000001000000101000", -- 4135 FREE #<CONS 0 4136>
 "00000000000000000001000000101001", -- 4136 FREE #<CONS 0 4137>
 "00000000000000000001000000101010", -- 4137 FREE #<CONS 0 4138>
 "00000000000000000001000000101011", -- 4138 FREE #<CONS 0 4139>
 "00000000000000000001000000101100", -- 4139 FREE #<CONS 0 4140>
 "00000000000000000001000000101101", -- 4140 FREE #<CONS 0 4141>
 "00000000000000000001000000101110", -- 4141 FREE #<CONS 0 4142>
 "00000000000000000001000000101111", -- 4142 FREE #<CONS 0 4143>
 "00000000000000000001000000110000", -- 4143 FREE #<CONS 0 4144>
 "00000000000000000001000000110001", -- 4144 FREE #<CONS 0 4145>
 "00000000000000000001000000110010", -- 4145 FREE #<CONS 0 4146>
 "00000000000000000001000000110011", -- 4146 FREE #<CONS 0 4147>
 "00000000000000000001000000110100", -- 4147 FREE #<CONS 0 4148>
 "00000000000000000001000000110101", -- 4148 FREE #<CONS 0 4149>
 "00000000000000000001000000110110", -- 4149 FREE #<CONS 0 4150>
 "00000000000000000001000000110111", -- 4150 FREE #<CONS 0 4151>
 "00000000000000000001000000111000", -- 4151 FREE #<CONS 0 4152>
 "00000000000000000001000000111001", -- 4152 FREE #<CONS 0 4153>
 "00000000000000000001000000111010", -- 4153 FREE #<CONS 0 4154>
 "00000000000000000001000000111011", -- 4154 FREE #<CONS 0 4155>
 "00000000000000000001000000111100", -- 4155 FREE #<CONS 0 4156>
 "00000000000000000001000000111101", -- 4156 FREE #<CONS 0 4157>
 "00000000000000000001000000111110", -- 4157 FREE #<CONS 0 4158>
 "00000000000000000001000000111111", -- 4158 FREE #<CONS 0 4159>
 "00000000000000000001000001000000", -- 4159 FREE #<CONS 0 4160>
 "00000000000000000001000001000001", -- 4160 FREE #<CONS 0 4161>
 "00000000000000000001000001000010", -- 4161 FREE #<CONS 0 4162>
 "00000000000000000001000001000011", -- 4162 FREE #<CONS 0 4163>
 "00000000000000000001000001000100", -- 4163 FREE #<CONS 0 4164>
 "00000000000000000001000001000101", -- 4164 FREE #<CONS 0 4165>
 "00000000000000000001000001000110", -- 4165 FREE #<CONS 0 4166>
 "00000000000000000001000001000111", -- 4166 FREE #<CONS 0 4167>
 "00000000000000000001000001001000", -- 4167 FREE #<CONS 0 4168>
 "00000000000000000001000001001001", -- 4168 FREE #<CONS 0 4169>
 "00000000000000000001000001001010", -- 4169 FREE #<CONS 0 4170>
 "00000000000000000001000001001011", -- 4170 FREE #<CONS 0 4171>
 "00000000000000000001000001001100", -- 4171 FREE #<CONS 0 4172>
 "00000000000000000001000001001101", -- 4172 FREE #<CONS 0 4173>
 "00000000000000000001000001001110", -- 4173 FREE #<CONS 0 4174>
 "00000000000000000001000001001111", -- 4174 FREE #<CONS 0 4175>
 "00000000000000000001000001010000", -- 4175 FREE #<CONS 0 4176>
 "00000000000000000001000001010001", -- 4176 FREE #<CONS 0 4177>
 "00000000000000000001000001010010", -- 4177 FREE #<CONS 0 4178>
 "00000000000000000001000001010011", -- 4178 FREE #<CONS 0 4179>
 "00000000000000000001000001010100", -- 4179 FREE #<CONS 0 4180>
 "00000000000000000001000001010101", -- 4180 FREE #<CONS 0 4181>
 "00000000000000000001000001010110", -- 4181 FREE #<CONS 0 4182>
 "00000000000000000001000001010111", -- 4182 FREE #<CONS 0 4183>
 "00000000000000000001000001011000", -- 4183 FREE #<CONS 0 4184>
 "00000000000000000001000001011001", -- 4184 FREE #<CONS 0 4185>
 "00000000000000000001000001011010", -- 4185 FREE #<CONS 0 4186>
 "00000000000000000001000001011011", -- 4186 FREE #<CONS 0 4187>
 "00000000000000000001000001011100", -- 4187 FREE #<CONS 0 4188>
 "00000000000000000001000001011101", -- 4188 FREE #<CONS 0 4189>
 "00000000000000000001000001011110", -- 4189 FREE #<CONS 0 4190>
 "00000000000000000001000001011111", -- 4190 FREE #<CONS 0 4191>
 "00000000000000000001000001100000", -- 4191 FREE #<CONS 0 4192>
 "00000000000000000001000001100001", -- 4192 FREE #<CONS 0 4193>
 "00000000000000000001000001100010", -- 4193 FREE #<CONS 0 4194>
 "00000000000000000001000001100011", -- 4194 FREE #<CONS 0 4195>
 "00000000000000000001000001100100", -- 4195 FREE #<CONS 0 4196>
 "00000000000000000001000001100101", -- 4196 FREE #<CONS 0 4197>
 "00000000000000000001000001100110", -- 4197 FREE #<CONS 0 4198>
 "00000000000000000001000001100111", -- 4198 FREE #<CONS 0 4199>
 "00000000000000000001000001101000", -- 4199 FREE #<CONS 0 4200>
 "00000000000000000001000001101001", -- 4200 FREE #<CONS 0 4201>
 "00000000000000000001000001101010", -- 4201 FREE #<CONS 0 4202>
 "00000000000000000001000001101011", -- 4202 FREE #<CONS 0 4203>
 "00000000000000000001000001101100", -- 4203 FREE #<CONS 0 4204>
 "00000000000000000001000001101101", -- 4204 FREE #<CONS 0 4205>
 "00000000000000000001000001101110", -- 4205 FREE #<CONS 0 4206>
 "00000000000000000001000001101111", -- 4206 FREE #<CONS 0 4207>
 "00000000000000000001000001110000", -- 4207 FREE #<CONS 0 4208>
 "00000000000000000001000001110001", -- 4208 FREE #<CONS 0 4209>
 "00000000000000000001000001110010", -- 4209 FREE #<CONS 0 4210>
 "00000000000000000001000001110011", -- 4210 FREE #<CONS 0 4211>
 "00000000000000000001000001110100", -- 4211 FREE #<CONS 0 4212>
 "00000000000000000001000001110101", -- 4212 FREE #<CONS 0 4213>
 "00000000000000000001000001110110", -- 4213 FREE #<CONS 0 4214>
 "00000000000000000001000001110111", -- 4214 FREE #<CONS 0 4215>
 "00000000000000000001000001111000", -- 4215 FREE #<CONS 0 4216>
 "00000000000000000001000001111001", -- 4216 FREE #<CONS 0 4217>
 "00000000000000000001000001111010", -- 4217 FREE #<CONS 0 4218>
 "00000000000000000001000001111011", -- 4218 FREE #<CONS 0 4219>
 "00000000000000000001000001111100", -- 4219 FREE #<CONS 0 4220>
 "00000000000000000001000001111101", -- 4220 FREE #<CONS 0 4221>
 "00000000000000000001000001111110", -- 4221 FREE #<CONS 0 4222>
 "00000000000000000001000001111111", -- 4222 FREE #<CONS 0 4223>
 "00000000000000000001000010000000", -- 4223 FREE #<CONS 0 4224>
 "00000000000000000001000010000001", -- 4224 FREE #<CONS 0 4225>
 "00000000000000000001000010000010", -- 4225 FREE #<CONS 0 4226>
 "00000000000000000001000010000011", -- 4226 FREE #<CONS 0 4227>
 "00000000000000000001000010000100", -- 4227 FREE #<CONS 0 4228>
 "00000000000000000001000010000101", -- 4228 FREE #<CONS 0 4229>
 "00000000000000000001000010000110", -- 4229 FREE #<CONS 0 4230>
 "00000000000000000001000010000111", -- 4230 FREE #<CONS 0 4231>
 "00000000000000000001000010001000", -- 4231 FREE #<CONS 0 4232>
 "00000000000000000001000010001001", -- 4232 FREE #<CONS 0 4233>
 "00000000000000000001000010001010", -- 4233 FREE #<CONS 0 4234>
 "00000000000000000001000010001011", -- 4234 FREE #<CONS 0 4235>
 "00000000000000000001000010001100", -- 4235 FREE #<CONS 0 4236>
 "00000000000000000001000010001101", -- 4236 FREE #<CONS 0 4237>
 "00000000000000000001000010001110", -- 4237 FREE #<CONS 0 4238>
 "00000000000000000001000010001111", -- 4238 FREE #<CONS 0 4239>
 "00000000000000000001000010010000", -- 4239 FREE #<CONS 0 4240>
 "00000000000000000001000010010001", -- 4240 FREE #<CONS 0 4241>
 "00000000000000000001000010010010", -- 4241 FREE #<CONS 0 4242>
 "00000000000000000001000010010011", -- 4242 FREE #<CONS 0 4243>
 "00000000000000000001000010010100", -- 4243 FREE #<CONS 0 4244>
 "00000000000000000001000010010101", -- 4244 FREE #<CONS 0 4245>
 "00000000000000000001000010010110", -- 4245 FREE #<CONS 0 4246>
 "00000000000000000001000010010111", -- 4246 FREE #<CONS 0 4247>
 "00000000000000000001000010011000", -- 4247 FREE #<CONS 0 4248>
 "00000000000000000001000010011001", -- 4248 FREE #<CONS 0 4249>
 "00000000000000000001000010011010", -- 4249 FREE #<CONS 0 4250>
 "00000000000000000001000010011011", -- 4250 FREE #<CONS 0 4251>
 "00000000000000000001000010011100", -- 4251 FREE #<CONS 0 4252>
 "00000000000000000001000010011101", -- 4252 FREE #<CONS 0 4253>
 "00000000000000000001000010011110", -- 4253 FREE #<CONS 0 4254>
 "00000000000000000001000010011111", -- 4254 FREE #<CONS 0 4255>
 "00000000000000000001000010100000", -- 4255 FREE #<CONS 0 4256>
 "00000000000000000001000010100001", -- 4256 FREE #<CONS 0 4257>
 "00000000000000000001000010100010", -- 4257 FREE #<CONS 0 4258>
 "00000000000000000001000010100011", -- 4258 FREE #<CONS 0 4259>
 "00000000000000000001000010100100", -- 4259 FREE #<CONS 0 4260>
 "00000000000000000001000010100101", -- 4260 FREE #<CONS 0 4261>
 "00000000000000000001000010100110", -- 4261 FREE #<CONS 0 4262>
 "00000000000000000001000010100111", -- 4262 FREE #<CONS 0 4263>
 "00000000000000000001000010101000", -- 4263 FREE #<CONS 0 4264>
 "00000000000000000001000010101001", -- 4264 FREE #<CONS 0 4265>
 "00000000000000000001000010101010", -- 4265 FREE #<CONS 0 4266>
 "00000000000000000001000010101011", -- 4266 FREE #<CONS 0 4267>
 "00000000000000000001000010101100", -- 4267 FREE #<CONS 0 4268>
 "00000000000000000001000010101101", -- 4268 FREE #<CONS 0 4269>
 "00000000000000000001000010101110", -- 4269 FREE #<CONS 0 4270>
 "00000000000000000001000010101111", -- 4270 FREE #<CONS 0 4271>
 "00000000000000000001000010110000", -- 4271 FREE #<CONS 0 4272>
 "00000000000000000001000010110001", -- 4272 FREE #<CONS 0 4273>
 "00000000000000000001000010110010", -- 4273 FREE #<CONS 0 4274>
 "00000000000000000001000010110011", -- 4274 FREE #<CONS 0 4275>
 "00000000000000000001000010110100", -- 4275 FREE #<CONS 0 4276>
 "00000000000000000001000010110101", -- 4276 FREE #<CONS 0 4277>
 "00000000000000000001000010110110", -- 4277 FREE #<CONS 0 4278>
 "00000000000000000001000010110111", -- 4278 FREE #<CONS 0 4279>
 "00000000000000000001000010111000", -- 4279 FREE #<CONS 0 4280>
 "00000000000000000001000010111001", -- 4280 FREE #<CONS 0 4281>
 "00000000000000000001000010111010", -- 4281 FREE #<CONS 0 4282>
 "00000000000000000001000010111011", -- 4282 FREE #<CONS 0 4283>
 "00000000000000000001000010111100", -- 4283 FREE #<CONS 0 4284>
 "00000000000000000001000010111101", -- 4284 FREE #<CONS 0 4285>
 "00000000000000000001000010111110", -- 4285 FREE #<CONS 0 4286>
 "00000000000000000001000010111111", -- 4286 FREE #<CONS 0 4287>
 "00000000000000000001000011000000", -- 4287 FREE #<CONS 0 4288>
 "00000000000000000001000011000001", -- 4288 FREE #<CONS 0 4289>
 "00000000000000000001000011000010", -- 4289 FREE #<CONS 0 4290>
 "00000000000000000001000011000011", -- 4290 FREE #<CONS 0 4291>
 "00000000000000000001000011000100", -- 4291 FREE #<CONS 0 4292>
 "00000000000000000001000011000101", -- 4292 FREE #<CONS 0 4293>
 "00000000000000000001000011000110", -- 4293 FREE #<CONS 0 4294>
 "00000000000000000001000011000111", -- 4294 FREE #<CONS 0 4295>
 "00000000000000000001000011001000", -- 4295 FREE #<CONS 0 4296>
 "00000000000000000001000011001001", -- 4296 FREE #<CONS 0 4297>
 "00000000000000000001000011001010", -- 4297 FREE #<CONS 0 4298>
 "00000000000000000001000011001011", -- 4298 FREE #<CONS 0 4299>
 "00000000000000000001000011001100", -- 4299 FREE #<CONS 0 4300>
 "00000000000000000001000011001101", -- 4300 FREE #<CONS 0 4301>
 "00000000000000000001000011001110", -- 4301 FREE #<CONS 0 4302>
 "00000000000000000001000011001111", -- 4302 FREE #<CONS 0 4303>
 "00000000000000000001000011010000", -- 4303 FREE #<CONS 0 4304>
 "00000000000000000001000011010001", -- 4304 FREE #<CONS 0 4305>
 "00000000000000000001000011010010", -- 4305 FREE #<CONS 0 4306>
 "00000000000000000001000011010011", -- 4306 FREE #<CONS 0 4307>
 "00000000000000000001000011010100", -- 4307 FREE #<CONS 0 4308>
 "00000000000000000001000011010101", -- 4308 FREE #<CONS 0 4309>
 "00000000000000000001000011010110", -- 4309 FREE #<CONS 0 4310>
 "00000000000000000001000011010111", -- 4310 FREE #<CONS 0 4311>
 "00000000000000000001000011011000", -- 4311 FREE #<CONS 0 4312>
 "00000000000000000001000011011001", -- 4312 FREE #<CONS 0 4313>
 "00000000000000000001000011011010", -- 4313 FREE #<CONS 0 4314>
 "00000000000000000001000011011011", -- 4314 FREE #<CONS 0 4315>
 "00000000000000000001000011011100", -- 4315 FREE #<CONS 0 4316>
 "00000000000000000001000011011101", -- 4316 FREE #<CONS 0 4317>
 "00000000000000000001000011011110", -- 4317 FREE #<CONS 0 4318>
 "00000000000000000001000011011111", -- 4318 FREE #<CONS 0 4319>
 "00000000000000000001000011100000", -- 4319 FREE #<CONS 0 4320>
 "00000000000000000001000011100001", -- 4320 FREE #<CONS 0 4321>
 "00000000000000000001000011100010", -- 4321 FREE #<CONS 0 4322>
 "00000000000000000001000011100011", -- 4322 FREE #<CONS 0 4323>
 "00000000000000000001000011100100", -- 4323 FREE #<CONS 0 4324>
 "00000000000000000001000011100101", -- 4324 FREE #<CONS 0 4325>
 "00000000000000000001000011100110", -- 4325 FREE #<CONS 0 4326>
 "00000000000000000001000011100111", -- 4326 FREE #<CONS 0 4327>
 "00000000000000000001000011101000", -- 4327 FREE #<CONS 0 4328>
 "00000000000000000001000011101001", -- 4328 FREE #<CONS 0 4329>
 "00000000000000000001000011101010", -- 4329 FREE #<CONS 0 4330>
 "00000000000000000001000011101011", -- 4330 FREE #<CONS 0 4331>
 "00000000000000000001000011101100", -- 4331 FREE #<CONS 0 4332>
 "00000000000000000001000011101101", -- 4332 FREE #<CONS 0 4333>
 "00000000000000000001000011101110", -- 4333 FREE #<CONS 0 4334>
 "00000000000000000001000011101111", -- 4334 FREE #<CONS 0 4335>
 "00000000000000000001000011110000", -- 4335 FREE #<CONS 0 4336>
 "00000000000000000001000011110001", -- 4336 FREE #<CONS 0 4337>
 "00000000000000000001000011110010", -- 4337 FREE #<CONS 0 4338>
 "00000000000000000001000011110011", -- 4338 FREE #<CONS 0 4339>
 "00000000000000000001000011110100", -- 4339 FREE #<CONS 0 4340>
 "00000000000000000001000011110101", -- 4340 FREE #<CONS 0 4341>
 "00000000000000000001000011110110", -- 4341 FREE #<CONS 0 4342>
 "00000000000000000001000011110111", -- 4342 FREE #<CONS 0 4343>
 "00000000000000000001000011111000", -- 4343 FREE #<CONS 0 4344>
 "00000000000000000001000011111001", -- 4344 FREE #<CONS 0 4345>
 "00000000000000000001000011111010", -- 4345 FREE #<CONS 0 4346>
 "00000000000000000001000011111011", -- 4346 FREE #<CONS 0 4347>
 "00000000000000000001000011111100", -- 4347 FREE #<CONS 0 4348>
 "00000000000000000001000011111101", -- 4348 FREE #<CONS 0 4349>
 "00000000000000000001000011111110", -- 4349 FREE #<CONS 0 4350>
 "00000000000000000001000011111111", -- 4350 FREE #<CONS 0 4351>
 "00000000000000000001000100000000", -- 4351 FREE #<CONS 0 4352>
 "00000000000000000001000100000001", -- 4352 FREE #<CONS 0 4353>
 "00000000000000000001000100000010", -- 4353 FREE #<CONS 0 4354>
 "00000000000000000001000100000011", -- 4354 FREE #<CONS 0 4355>
 "00000000000000000001000100000100", -- 4355 FREE #<CONS 0 4356>
 "00000000000000000001000100000101", -- 4356 FREE #<CONS 0 4357>
 "00000000000000000001000100000110", -- 4357 FREE #<CONS 0 4358>
 "00000000000000000001000100000111", -- 4358 FREE #<CONS 0 4359>
 "00000000000000000001000100001000", -- 4359 FREE #<CONS 0 4360>
 "00000000000000000001000100001001", -- 4360 FREE #<CONS 0 4361>
 "00000000000000000001000100001010", -- 4361 FREE #<CONS 0 4362>
 "00000000000000000001000100001011", -- 4362 FREE #<CONS 0 4363>
 "00000000000000000001000100001100", -- 4363 FREE #<CONS 0 4364>
 "00000000000000000001000100001101", -- 4364 FREE #<CONS 0 4365>
 "00000000000000000001000100001110", -- 4365 FREE #<CONS 0 4366>
 "00000000000000000001000100001111", -- 4366 FREE #<CONS 0 4367>
 "00000000000000000001000100010000", -- 4367 FREE #<CONS 0 4368>
 "00000000000000000001000100010001", -- 4368 FREE #<CONS 0 4369>
 "00000000000000000001000100010010", -- 4369 FREE #<CONS 0 4370>
 "00000000000000000001000100010011", -- 4370 FREE #<CONS 0 4371>
 "00000000000000000001000100010100", -- 4371 FREE #<CONS 0 4372>
 "00000000000000000001000100010101", -- 4372 FREE #<CONS 0 4373>
 "00000000000000000001000100010110", -- 4373 FREE #<CONS 0 4374>
 "00000000000000000001000100010111", -- 4374 FREE #<CONS 0 4375>
 "00000000000000000001000100011000", -- 4375 FREE #<CONS 0 4376>
 "00000000000000000001000100011001", -- 4376 FREE #<CONS 0 4377>
 "00000000000000000001000100011010", -- 4377 FREE #<CONS 0 4378>
 "00000000000000000001000100011011", -- 4378 FREE #<CONS 0 4379>
 "00000000000000000001000100011100", -- 4379 FREE #<CONS 0 4380>
 "00000000000000000001000100011101", -- 4380 FREE #<CONS 0 4381>
 "00000000000000000001000100011110", -- 4381 FREE #<CONS 0 4382>
 "00000000000000000001000100011111", -- 4382 FREE #<CONS 0 4383>
 "00000000000000000001000100100000", -- 4383 FREE #<CONS 0 4384>
 "00000000000000000001000100100001", -- 4384 FREE #<CONS 0 4385>
 "00000000000000000001000100100010", -- 4385 FREE #<CONS 0 4386>
 "00000000000000000001000100100011", -- 4386 FREE #<CONS 0 4387>
 "00000000000000000001000100100100", -- 4387 FREE #<CONS 0 4388>
 "00000000000000000001000100100101", -- 4388 FREE #<CONS 0 4389>
 "00000000000000000001000100100110", -- 4389 FREE #<CONS 0 4390>
 "00000000000000000001000100100111", -- 4390 FREE #<CONS 0 4391>
 "00000000000000000001000100101000", -- 4391 FREE #<CONS 0 4392>
 "00000000000000000001000100101001", -- 4392 FREE #<CONS 0 4393>
 "00000000000000000001000100101010", -- 4393 FREE #<CONS 0 4394>
 "00000000000000000001000100101011", -- 4394 FREE #<CONS 0 4395>
 "00000000000000000001000100101100", -- 4395 FREE #<CONS 0 4396>
 "00000000000000000001000100101101", -- 4396 FREE #<CONS 0 4397>
 "00000000000000000001000100101110", -- 4397 FREE #<CONS 0 4398>
 "00000000000000000001000100101111", -- 4398 FREE #<CONS 0 4399>
 "00000000000000000001000100110000", -- 4399 FREE #<CONS 0 4400>
 "00000000000000000001000100110001", -- 4400 FREE #<CONS 0 4401>
 "00000000000000000001000100110010", -- 4401 FREE #<CONS 0 4402>
 "00000000000000000001000100110011", -- 4402 FREE #<CONS 0 4403>
 "00000000000000000001000100110100", -- 4403 FREE #<CONS 0 4404>
 "00000000000000000001000100110101", -- 4404 FREE #<CONS 0 4405>
 "00000000000000000001000100110110", -- 4405 FREE #<CONS 0 4406>
 "00000000000000000001000100110111", -- 4406 FREE #<CONS 0 4407>
 "00000000000000000001000100111000", -- 4407 FREE #<CONS 0 4408>
 "00000000000000000001000100111001", -- 4408 FREE #<CONS 0 4409>
 "00000000000000000001000100111010", -- 4409 FREE #<CONS 0 4410>
 "00000000000000000001000100111011", -- 4410 FREE #<CONS 0 4411>
 "00000000000000000001000100111100", -- 4411 FREE #<CONS 0 4412>
 "00000000000000000001000100111101", -- 4412 FREE #<CONS 0 4413>
 "00000000000000000001000100111110", -- 4413 FREE #<CONS 0 4414>
 "00000000000000000001000100111111", -- 4414 FREE #<CONS 0 4415>
 "00000000000000000001000101000000", -- 4415 FREE #<CONS 0 4416>
 "00000000000000000001000101000001", -- 4416 FREE #<CONS 0 4417>
 "00000000000000000001000101000010", -- 4417 FREE #<CONS 0 4418>
 "00000000000000000001000101000011", -- 4418 FREE #<CONS 0 4419>
 "00000000000000000001000101000100", -- 4419 FREE #<CONS 0 4420>
 "00000000000000000001000101000101", -- 4420 FREE #<CONS 0 4421>
 "00000000000000000001000101000110", -- 4421 FREE #<CONS 0 4422>
 "00000000000000000001000101000111", -- 4422 FREE #<CONS 0 4423>
 "00000000000000000001000101001000", -- 4423 FREE #<CONS 0 4424>
 "00000000000000000001000101001001", -- 4424 FREE #<CONS 0 4425>
 "00000000000000000001000101001010", -- 4425 FREE #<CONS 0 4426>
 "00000000000000000001000101001011", -- 4426 FREE #<CONS 0 4427>
 "00000000000000000001000101001100", -- 4427 FREE #<CONS 0 4428>
 "00000000000000000001000101001101", -- 4428 FREE #<CONS 0 4429>
 "00000000000000000001000101001110", -- 4429 FREE #<CONS 0 4430>
 "00000000000000000001000101001111", -- 4430 FREE #<CONS 0 4431>
 "00000000000000000001000101010000", -- 4431 FREE #<CONS 0 4432>
 "00000000000000000001000101010001", -- 4432 FREE #<CONS 0 4433>
 "00000000000000000001000101010010", -- 4433 FREE #<CONS 0 4434>
 "00000000000000000001000101010011", -- 4434 FREE #<CONS 0 4435>
 "00000000000000000001000101010100", -- 4435 FREE #<CONS 0 4436>
 "00000000000000000001000101010101", -- 4436 FREE #<CONS 0 4437>
 "00000000000000000001000101010110", -- 4437 FREE #<CONS 0 4438>
 "00000000000000000001000101010111", -- 4438 FREE #<CONS 0 4439>
 "00000000000000000001000101011000", -- 4439 FREE #<CONS 0 4440>
 "00000000000000000001000101011001", -- 4440 FREE #<CONS 0 4441>
 "00000000000000000001000101011010", -- 4441 FREE #<CONS 0 4442>
 "00000000000000000001000101011011", -- 4442 FREE #<CONS 0 4443>
 "00000000000000000001000101011100", -- 4443 FREE #<CONS 0 4444>
 "00000000000000000001000101011101", -- 4444 FREE #<CONS 0 4445>
 "00000000000000000001000101011110", -- 4445 FREE #<CONS 0 4446>
 "00000000000000000001000101011111", -- 4446 FREE #<CONS 0 4447>
 "00000000000000000001000101100000", -- 4447 FREE #<CONS 0 4448>
 "00000000000000000001000101100001", -- 4448 FREE #<CONS 0 4449>
 "00000000000000000001000101100010", -- 4449 FREE #<CONS 0 4450>
 "00000000000000000001000101100011", -- 4450 FREE #<CONS 0 4451>
 "00000000000000000001000101100100", -- 4451 FREE #<CONS 0 4452>
 "00000000000000000001000101100101", -- 4452 FREE #<CONS 0 4453>
 "00000000000000000001000101100110", -- 4453 FREE #<CONS 0 4454>
 "00000000000000000001000101100111", -- 4454 FREE #<CONS 0 4455>
 "00000000000000000001000101101000", -- 4455 FREE #<CONS 0 4456>
 "00000000000000000001000101101001", -- 4456 FREE #<CONS 0 4457>
 "00000000000000000001000101101010", -- 4457 FREE #<CONS 0 4458>
 "00000000000000000001000101101011", -- 4458 FREE #<CONS 0 4459>
 "00000000000000000001000101101100", -- 4459 FREE #<CONS 0 4460>
 "00000000000000000001000101101101", -- 4460 FREE #<CONS 0 4461>
 "00000000000000000001000101101110", -- 4461 FREE #<CONS 0 4462>
 "00000000000000000001000101101111", -- 4462 FREE #<CONS 0 4463>
 "00000000000000000001000101110000", -- 4463 FREE #<CONS 0 4464>
 "00000000000000000001000101110001", -- 4464 FREE #<CONS 0 4465>
 "00000000000000000001000101110010", -- 4465 FREE #<CONS 0 4466>
 "00000000000000000001000101110011", -- 4466 FREE #<CONS 0 4467>
 "00000000000000000001000101110100", -- 4467 FREE #<CONS 0 4468>
 "00000000000000000001000101110101", -- 4468 FREE #<CONS 0 4469>
 "00000000000000000001000101110110", -- 4469 FREE #<CONS 0 4470>
 "00000000000000000001000101110111", -- 4470 FREE #<CONS 0 4471>
 "00000000000000000001000101111000", -- 4471 FREE #<CONS 0 4472>
 "00000000000000000001000101111001", -- 4472 FREE #<CONS 0 4473>
 "00000000000000000001000101111010", -- 4473 FREE #<CONS 0 4474>
 "00000000000000000001000101111011", -- 4474 FREE #<CONS 0 4475>
 "00000000000000000001000101111100", -- 4475 FREE #<CONS 0 4476>
 "00000000000000000001000101111101", -- 4476 FREE #<CONS 0 4477>
 "00000000000000000001000101111110", -- 4477 FREE #<CONS 0 4478>
 "00000000000000000001000101111111", -- 4478 FREE #<CONS 0 4479>
 "00000000000000000001000110000000", -- 4479 FREE #<CONS 0 4480>
 "00000000000000000001000110000001", -- 4480 FREE #<CONS 0 4481>
 "00000000000000000001000110000010", -- 4481 FREE #<CONS 0 4482>
 "00000000000000000001000110000011", -- 4482 FREE #<CONS 0 4483>
 "00000000000000000001000110000100", -- 4483 FREE #<CONS 0 4484>
 "00000000000000000001000110000101", -- 4484 FREE #<CONS 0 4485>
 "00000000000000000001000110000110", -- 4485 FREE #<CONS 0 4486>
 "00000000000000000001000110000111", -- 4486 FREE #<CONS 0 4487>
 "00000000000000000001000110001000", -- 4487 FREE #<CONS 0 4488>
 "00000000000000000001000110001001", -- 4488 FREE #<CONS 0 4489>
 "00000000000000000001000110001010", -- 4489 FREE #<CONS 0 4490>
 "00000000000000000001000110001011", -- 4490 FREE #<CONS 0 4491>
 "00000000000000000001000110001100", -- 4491 FREE #<CONS 0 4492>
 "00000000000000000001000110001101", -- 4492 FREE #<CONS 0 4493>
 "00000000000000000001000110001110", -- 4493 FREE #<CONS 0 4494>
 "00000000000000000001000110001111", -- 4494 FREE #<CONS 0 4495>
 "00000000000000000001000110010000", -- 4495 FREE #<CONS 0 4496>
 "00000000000000000001000110010001", -- 4496 FREE #<CONS 0 4497>
 "00000000000000000001000110010010", -- 4497 FREE #<CONS 0 4498>
 "00000000000000000001000110010011", -- 4498 FREE #<CONS 0 4499>
 "00000000000000000001000110010100", -- 4499 FREE #<CONS 0 4500>
 "00000000000000000001000110010101", -- 4500 FREE #<CONS 0 4501>
 "00000000000000000001000110010110", -- 4501 FREE #<CONS 0 4502>
 "00000000000000000001000110010111", -- 4502 FREE #<CONS 0 4503>
 "00000000000000000001000110011000", -- 4503 FREE #<CONS 0 4504>
 "00000000000000000001000110011001", -- 4504 FREE #<CONS 0 4505>
 "00000000000000000001000110011010", -- 4505 FREE #<CONS 0 4506>
 "00000000000000000001000110011011", -- 4506 FREE #<CONS 0 4507>
 "00000000000000000001000110011100", -- 4507 FREE #<CONS 0 4508>
 "00000000000000000001000110011101", -- 4508 FREE #<CONS 0 4509>
 "00000000000000000001000110011110", -- 4509 FREE #<CONS 0 4510>
 "00000000000000000001000110011111", -- 4510 FREE #<CONS 0 4511>
 "00000000000000000001000110100000", -- 4511 FREE #<CONS 0 4512>
 "00000000000000000001000110100001", -- 4512 FREE #<CONS 0 4513>
 "00000000000000000001000110100010", -- 4513 FREE #<CONS 0 4514>
 "00000000000000000001000110100011", -- 4514 FREE #<CONS 0 4515>
 "00000000000000000001000110100100", -- 4515 FREE #<CONS 0 4516>
 "00000000000000000001000110100101", -- 4516 FREE #<CONS 0 4517>
 "00000000000000000001000110100110", -- 4517 FREE #<CONS 0 4518>
 "00000000000000000001000110100111", -- 4518 FREE #<CONS 0 4519>
 "00000000000000000001000110101000", -- 4519 FREE #<CONS 0 4520>
 "00000000000000000001000110101001", -- 4520 FREE #<CONS 0 4521>
 "00000000000000000001000110101010", -- 4521 FREE #<CONS 0 4522>
 "00000000000000000001000110101011", -- 4522 FREE #<CONS 0 4523>
 "00000000000000000001000110101100", -- 4523 FREE #<CONS 0 4524>
 "00000000000000000001000110101101", -- 4524 FREE #<CONS 0 4525>
 "00000000000000000001000110101110", -- 4525 FREE #<CONS 0 4526>
 "00000000000000000001000110101111", -- 4526 FREE #<CONS 0 4527>
 "00000000000000000001000110110000", -- 4527 FREE #<CONS 0 4528>
 "00000000000000000001000110110001", -- 4528 FREE #<CONS 0 4529>
 "00000000000000000001000110110010", -- 4529 FREE #<CONS 0 4530>
 "00000000000000000001000110110011", -- 4530 FREE #<CONS 0 4531>
 "00000000000000000001000110110100", -- 4531 FREE #<CONS 0 4532>
 "00000000000000000001000110110101", -- 4532 FREE #<CONS 0 4533>
 "00000000000000000001000110110110", -- 4533 FREE #<CONS 0 4534>
 "00000000000000000001000110110111", -- 4534 FREE #<CONS 0 4535>
 "00000000000000000001000110111000", -- 4535 FREE #<CONS 0 4536>
 "00000000000000000001000110111001", -- 4536 FREE #<CONS 0 4537>
 "00000000000000000001000110111010", -- 4537 FREE #<CONS 0 4538>
 "00000000000000000001000110111011", -- 4538 FREE #<CONS 0 4539>
 "00000000000000000001000110111100", -- 4539 FREE #<CONS 0 4540>
 "00000000000000000001000110111101", -- 4540 FREE #<CONS 0 4541>
 "00000000000000000001000110111110", -- 4541 FREE #<CONS 0 4542>
 "00000000000000000001000110111111", -- 4542 FREE #<CONS 0 4543>
 "00000000000000000001000111000000", -- 4543 FREE #<CONS 0 4544>
 "00000000000000000001000111000001", -- 4544 FREE #<CONS 0 4545>
 "00000000000000000001000111000010", -- 4545 FREE #<CONS 0 4546>
 "00000000000000000001000111000011", -- 4546 FREE #<CONS 0 4547>
 "00000000000000000001000111000100", -- 4547 FREE #<CONS 0 4548>
 "00000000000000000001000111000101", -- 4548 FREE #<CONS 0 4549>
 "00000000000000000001000111000110", -- 4549 FREE #<CONS 0 4550>
 "00000000000000000001000111000111", -- 4550 FREE #<CONS 0 4551>
 "00000000000000000001000111001000", -- 4551 FREE #<CONS 0 4552>
 "00000000000000000001000111001001", -- 4552 FREE #<CONS 0 4553>
 "00000000000000000001000111001010", -- 4553 FREE #<CONS 0 4554>
 "00000000000000000001000111001011", -- 4554 FREE #<CONS 0 4555>
 "00000000000000000001000111001100", -- 4555 FREE #<CONS 0 4556>
 "00000000000000000001000111001101", -- 4556 FREE #<CONS 0 4557>
 "00000000000000000001000111001110", -- 4557 FREE #<CONS 0 4558>
 "00000000000000000001000111001111", -- 4558 FREE #<CONS 0 4559>
 "00000000000000000001000111010000", -- 4559 FREE #<CONS 0 4560>
 "00000000000000000001000111010001", -- 4560 FREE #<CONS 0 4561>
 "00000000000000000001000111010010", -- 4561 FREE #<CONS 0 4562>
 "00000000000000000001000111010011", -- 4562 FREE #<CONS 0 4563>
 "00000000000000000001000111010100", -- 4563 FREE #<CONS 0 4564>
 "00000000000000000001000111010101", -- 4564 FREE #<CONS 0 4565>
 "00000000000000000001000111010110", -- 4565 FREE #<CONS 0 4566>
 "00000000000000000001000111010111", -- 4566 FREE #<CONS 0 4567>
 "00000000000000000001000111011000", -- 4567 FREE #<CONS 0 4568>
 "00000000000000000001000111011001", -- 4568 FREE #<CONS 0 4569>
 "00000000000000000001000111011010", -- 4569 FREE #<CONS 0 4570>
 "00000000000000000001000111011011", -- 4570 FREE #<CONS 0 4571>
 "00000000000000000001000111011100", -- 4571 FREE #<CONS 0 4572>
 "00000000000000000001000111011101", -- 4572 FREE #<CONS 0 4573>
 "00000000000000000001000111011110", -- 4573 FREE #<CONS 0 4574>
 "00000000000000000001000111011111", -- 4574 FREE #<CONS 0 4575>
 "00000000000000000001000111100000", -- 4575 FREE #<CONS 0 4576>
 "00000000000000000001000111100001", -- 4576 FREE #<CONS 0 4577>
 "00000000000000000001000111100010", -- 4577 FREE #<CONS 0 4578>
 "00000000000000000001000111100011", -- 4578 FREE #<CONS 0 4579>
 "00000000000000000001000111100100", -- 4579 FREE #<CONS 0 4580>
 "00000000000000000001000111100101", -- 4580 FREE #<CONS 0 4581>
 "00000000000000000001000111100110", -- 4581 FREE #<CONS 0 4582>
 "00000000000000000001000111100111", -- 4582 FREE #<CONS 0 4583>
 "00000000000000000001000111101000", -- 4583 FREE #<CONS 0 4584>
 "00000000000000000001000111101001", -- 4584 FREE #<CONS 0 4585>
 "00000000000000000001000111101010", -- 4585 FREE #<CONS 0 4586>
 "00000000000000000001000111101011", -- 4586 FREE #<CONS 0 4587>
 "00000000000000000001000111101100", -- 4587 FREE #<CONS 0 4588>
 "00000000000000000001000111101101", -- 4588 FREE #<CONS 0 4589>
 "00000000000000000001000111101110", -- 4589 FREE #<CONS 0 4590>
 "00000000000000000001000111101111", -- 4590 FREE #<CONS 0 4591>
 "00000000000000000001000111110000", -- 4591 FREE #<CONS 0 4592>
 "00000000000000000001000111110001", -- 4592 FREE #<CONS 0 4593>
 "00000000000000000001000111110010", -- 4593 FREE #<CONS 0 4594>
 "00000000000000000001000111110011", -- 4594 FREE #<CONS 0 4595>
 "00000000000000000001000111110100", -- 4595 FREE #<CONS 0 4596>
 "00000000000000000001000111110101", -- 4596 FREE #<CONS 0 4597>
 "00000000000000000001000111110110", -- 4597 FREE #<CONS 0 4598>
 "00000000000000000001000111110111", -- 4598 FREE #<CONS 0 4599>
 "00000000000000000001000111111000", -- 4599 FREE #<CONS 0 4600>
 "00000000000000000001000111111001", -- 4600 FREE #<CONS 0 4601>
 "00000000000000000001000111111010", -- 4601 FREE #<CONS 0 4602>
 "00000000000000000001000111111011", -- 4602 FREE #<CONS 0 4603>
 "00000000000000000001000111111100", -- 4603 FREE #<CONS 0 4604>
 "00000000000000000001000111111101", -- 4604 FREE #<CONS 0 4605>
 "00000000000000000001000111111110", -- 4605 FREE #<CONS 0 4606>
 "00000000000000000001000111111111", -- 4606 FREE #<CONS 0 4607>
 "00000000000000000001001000000000", -- 4607 FREE #<CONS 0 4608>
 "00000000000000000001001000000001", -- 4608 FREE #<CONS 0 4609>
 "00000000000000000001001000000010", -- 4609 FREE #<CONS 0 4610>
 "00000000000000000001001000000011", -- 4610 FREE #<CONS 0 4611>
 "00000000000000000001001000000100", -- 4611 FREE #<CONS 0 4612>
 "00000000000000000001001000000101", -- 4612 FREE #<CONS 0 4613>
 "00000000000000000001001000000110", -- 4613 FREE #<CONS 0 4614>
 "00000000000000000001001000000111", -- 4614 FREE #<CONS 0 4615>
 "00000000000000000001001000001000", -- 4615 FREE #<CONS 0 4616>
 "00000000000000000001001000001001", -- 4616 FREE #<CONS 0 4617>
 "00000000000000000001001000001010", -- 4617 FREE #<CONS 0 4618>
 "00000000000000000001001000001011", -- 4618 FREE #<CONS 0 4619>
 "00000000000000000001001000001100", -- 4619 FREE #<CONS 0 4620>
 "00000000000000000001001000001101", -- 4620 FREE #<CONS 0 4621>
 "00000000000000000001001000001110", -- 4621 FREE #<CONS 0 4622>
 "00000000000000000001001000001111", -- 4622 FREE #<CONS 0 4623>
 "00000000000000000001001000010000", -- 4623 FREE #<CONS 0 4624>
 "00000000000000000001001000010001", -- 4624 FREE #<CONS 0 4625>
 "00000000000000000001001000010010", -- 4625 FREE #<CONS 0 4626>
 "00000000000000000001001000010011", -- 4626 FREE #<CONS 0 4627>
 "00000000000000000001001000010100", -- 4627 FREE #<CONS 0 4628>
 "00000000000000000001001000010101", -- 4628 FREE #<CONS 0 4629>
 "00000000000000000001001000010110", -- 4629 FREE #<CONS 0 4630>
 "00000000000000000001001000010111", -- 4630 FREE #<CONS 0 4631>
 "00000000000000000001001000011000", -- 4631 FREE #<CONS 0 4632>
 "00000000000000000001001000011001", -- 4632 FREE #<CONS 0 4633>
 "00000000000000000001001000011010", -- 4633 FREE #<CONS 0 4634>
 "00000000000000000001001000011011", -- 4634 FREE #<CONS 0 4635>
 "00000000000000000001001000011100", -- 4635 FREE #<CONS 0 4636>
 "00000000000000000001001000011101", -- 4636 FREE #<CONS 0 4637>
 "00000000000000000001001000011110", -- 4637 FREE #<CONS 0 4638>
 "00000000000000000001001000011111", -- 4638 FREE #<CONS 0 4639>
 "00000000000000000001001000100000", -- 4639 FREE #<CONS 0 4640>
 "00000000000000000001001000100001", -- 4640 FREE #<CONS 0 4641>
 "00000000000000000001001000100010", -- 4641 FREE #<CONS 0 4642>
 "00000000000000000001001000100011", -- 4642 FREE #<CONS 0 4643>
 "00000000000000000001001000100100", -- 4643 FREE #<CONS 0 4644>
 "00000000000000000001001000100101", -- 4644 FREE #<CONS 0 4645>
 "00000000000000000001001000100110", -- 4645 FREE #<CONS 0 4646>
 "00000000000000000001001000100111", -- 4646 FREE #<CONS 0 4647>
 "00000000000000000001001000101000", -- 4647 FREE #<CONS 0 4648>
 "00000000000000000001001000101001", -- 4648 FREE #<CONS 0 4649>
 "00000000000000000001001000101010", -- 4649 FREE #<CONS 0 4650>
 "00000000000000000001001000101011", -- 4650 FREE #<CONS 0 4651>
 "00000000000000000001001000101100", -- 4651 FREE #<CONS 0 4652>
 "00000000000000000001001000101101", -- 4652 FREE #<CONS 0 4653>
 "00000000000000000001001000101110", -- 4653 FREE #<CONS 0 4654>
 "00000000000000000001001000101111", -- 4654 FREE #<CONS 0 4655>
 "00000000000000000001001000110000", -- 4655 FREE #<CONS 0 4656>
 "00000000000000000001001000110001", -- 4656 FREE #<CONS 0 4657>
 "00000000000000000001001000110010", -- 4657 FREE #<CONS 0 4658>
 "00000000000000000001001000110011", -- 4658 FREE #<CONS 0 4659>
 "00000000000000000001001000110100", -- 4659 FREE #<CONS 0 4660>
 "00000000000000000001001000110101", -- 4660 FREE #<CONS 0 4661>
 "00000000000000000001001000110110", -- 4661 FREE #<CONS 0 4662>
 "00000000000000000001001000110111", -- 4662 FREE #<CONS 0 4663>
 "00000000000000000001001000111000", -- 4663 FREE #<CONS 0 4664>
 "00000000000000000001001000111001", -- 4664 FREE #<CONS 0 4665>
 "00000000000000000001001000111010", -- 4665 FREE #<CONS 0 4666>
 "00000000000000000001001000111011", -- 4666 FREE #<CONS 0 4667>
 "00000000000000000001001000111100", -- 4667 FREE #<CONS 0 4668>
 "00000000000000000001001000111101", -- 4668 FREE #<CONS 0 4669>
 "00000000000000000001001000111110", -- 4669 FREE #<CONS 0 4670>
 "00000000000000000001001000111111", -- 4670 FREE #<CONS 0 4671>
 "00000000000000000001001001000000", -- 4671 FREE #<CONS 0 4672>
 "00000000000000000001001001000001", -- 4672 FREE #<CONS 0 4673>
 "00000000000000000001001001000010", -- 4673 FREE #<CONS 0 4674>
 "00000000000000000001001001000011", -- 4674 FREE #<CONS 0 4675>
 "00000000000000000001001001000100", -- 4675 FREE #<CONS 0 4676>
 "00000000000000000001001001000101", -- 4676 FREE #<CONS 0 4677>
 "00000000000000000001001001000110", -- 4677 FREE #<CONS 0 4678>
 "00000000000000000001001001000111", -- 4678 FREE #<CONS 0 4679>
 "00000000000000000001001001001000", -- 4679 FREE #<CONS 0 4680>
 "00000000000000000001001001001001", -- 4680 FREE #<CONS 0 4681>
 "00000000000000000001001001001010", -- 4681 FREE #<CONS 0 4682>
 "00000000000000000001001001001011", -- 4682 FREE #<CONS 0 4683>
 "00000000000000000001001001001100", -- 4683 FREE #<CONS 0 4684>
 "00000000000000000001001001001101", -- 4684 FREE #<CONS 0 4685>
 "00000000000000000001001001001110", -- 4685 FREE #<CONS 0 4686>
 "00000000000000000001001001001111", -- 4686 FREE #<CONS 0 4687>
 "00000000000000000001001001010000", -- 4687 FREE #<CONS 0 4688>
 "00000000000000000001001001010001", -- 4688 FREE #<CONS 0 4689>
 "00000000000000000001001001010010", -- 4689 FREE #<CONS 0 4690>
 "00000000000000000001001001010011", -- 4690 FREE #<CONS 0 4691>
 "00000000000000000001001001010100", -- 4691 FREE #<CONS 0 4692>
 "00000000000000000001001001010101", -- 4692 FREE #<CONS 0 4693>
 "00000000000000000001001001010110", -- 4693 FREE #<CONS 0 4694>
 "00000000000000000001001001010111", -- 4694 FREE #<CONS 0 4695>
 "00000000000000000001001001011000", -- 4695 FREE #<CONS 0 4696>
 "00000000000000000001001001011001", -- 4696 FREE #<CONS 0 4697>
 "00000000000000000001001001011010", -- 4697 FREE #<CONS 0 4698>
 "00000000000000000001001001011011", -- 4698 FREE #<CONS 0 4699>
 "00000000000000000001001001011100", -- 4699 FREE #<CONS 0 4700>
 "00000000000000000001001001011101", -- 4700 FREE #<CONS 0 4701>
 "00000000000000000001001001011110", -- 4701 FREE #<CONS 0 4702>
 "00000000000000000001001001011111", -- 4702 FREE #<CONS 0 4703>
 "00000000000000000001001001100000", -- 4703 FREE #<CONS 0 4704>
 "00000000000000000001001001100001", -- 4704 FREE #<CONS 0 4705>
 "00000000000000000001001001100010", -- 4705 FREE #<CONS 0 4706>
 "00000000000000000001001001100011", -- 4706 FREE #<CONS 0 4707>
 "00000000000000000001001001100100", -- 4707 FREE #<CONS 0 4708>
 "00000000000000000001001001100101", -- 4708 FREE #<CONS 0 4709>
 "00000000000000000001001001100110", -- 4709 FREE #<CONS 0 4710>
 "00000000000000000001001001100111", -- 4710 FREE #<CONS 0 4711>
 "00000000000000000001001001101000", -- 4711 FREE #<CONS 0 4712>
 "00000000000000000001001001101001", -- 4712 FREE #<CONS 0 4713>
 "00000000000000000001001001101010", -- 4713 FREE #<CONS 0 4714>
 "00000000000000000001001001101011", -- 4714 FREE #<CONS 0 4715>
 "00000000000000000001001001101100", -- 4715 FREE #<CONS 0 4716>
 "00000000000000000001001001101101", -- 4716 FREE #<CONS 0 4717>
 "00000000000000000001001001101110", -- 4717 FREE #<CONS 0 4718>
 "00000000000000000001001001101111", -- 4718 FREE #<CONS 0 4719>
 "00000000000000000001001001110000", -- 4719 FREE #<CONS 0 4720>
 "00000000000000000001001001110001", -- 4720 FREE #<CONS 0 4721>
 "00000000000000000001001001110010", -- 4721 FREE #<CONS 0 4722>
 "00000000000000000001001001110011", -- 4722 FREE #<CONS 0 4723>
 "00000000000000000001001001110100", -- 4723 FREE #<CONS 0 4724>
 "00000000000000000001001001110101", -- 4724 FREE #<CONS 0 4725>
 "00000000000000000001001001110110", -- 4725 FREE #<CONS 0 4726>
 "00000000000000000001001001110111", -- 4726 FREE #<CONS 0 4727>
 "00000000000000000001001001111000", -- 4727 FREE #<CONS 0 4728>
 "00000000000000000001001001111001", -- 4728 FREE #<CONS 0 4729>
 "00000000000000000001001001111010", -- 4729 FREE #<CONS 0 4730>
 "00000000000000000001001001111011", -- 4730 FREE #<CONS 0 4731>
 "00000000000000000001001001111100", -- 4731 FREE #<CONS 0 4732>
 "00000000000000000001001001111101", -- 4732 FREE #<CONS 0 4733>
 "00000000000000000001001001111110", -- 4733 FREE #<CONS 0 4734>
 "00000000000000000001001001111111", -- 4734 FREE #<CONS 0 4735>
 "00000000000000000001001010000000", -- 4735 FREE #<CONS 0 4736>
 "00000000000000000001001010000001", -- 4736 FREE #<CONS 0 4737>
 "00000000000000000001001010000010", -- 4737 FREE #<CONS 0 4738>
 "00000000000000000001001010000011", -- 4738 FREE #<CONS 0 4739>
 "00000000000000000001001010000100", -- 4739 FREE #<CONS 0 4740>
 "00000000000000000001001010000101", -- 4740 FREE #<CONS 0 4741>
 "00000000000000000001001010000110", -- 4741 FREE #<CONS 0 4742>
 "00000000000000000001001010000111", -- 4742 FREE #<CONS 0 4743>
 "00000000000000000001001010001000", -- 4743 FREE #<CONS 0 4744>
 "00000000000000000001001010001001", -- 4744 FREE #<CONS 0 4745>
 "00000000000000000001001010001010", -- 4745 FREE #<CONS 0 4746>
 "00000000000000000001001010001011", -- 4746 FREE #<CONS 0 4747>
 "00000000000000000001001010001100", -- 4747 FREE #<CONS 0 4748>
 "00000000000000000001001010001101", -- 4748 FREE #<CONS 0 4749>
 "00000000000000000001001010001110", -- 4749 FREE #<CONS 0 4750>
 "00000000000000000001001010001111", -- 4750 FREE #<CONS 0 4751>
 "00000000000000000001001010010000", -- 4751 FREE #<CONS 0 4752>
 "00000000000000000001001010010001", -- 4752 FREE #<CONS 0 4753>
 "00000000000000000001001010010010", -- 4753 FREE #<CONS 0 4754>
 "00000000000000000001001010010011", -- 4754 FREE #<CONS 0 4755>
 "00000000000000000001001010010100", -- 4755 FREE #<CONS 0 4756>
 "00000000000000000001001010010101", -- 4756 FREE #<CONS 0 4757>
 "00000000000000000001001010010110", -- 4757 FREE #<CONS 0 4758>
 "00000000000000000001001010010111", -- 4758 FREE #<CONS 0 4759>
 "00000000000000000001001010011000", -- 4759 FREE #<CONS 0 4760>
 "00000000000000000001001010011001", -- 4760 FREE #<CONS 0 4761>
 "00000000000000000001001010011010", -- 4761 FREE #<CONS 0 4762>
 "00000000000000000001001010011011", -- 4762 FREE #<CONS 0 4763>
 "00000000000000000001001010011100", -- 4763 FREE #<CONS 0 4764>
 "00000000000000000001001010011101", -- 4764 FREE #<CONS 0 4765>
 "00000000000000000001001010011110", -- 4765 FREE #<CONS 0 4766>
 "00000000000000000001001010011111", -- 4766 FREE #<CONS 0 4767>
 "00000000000000000001001010100000", -- 4767 FREE #<CONS 0 4768>
 "00000000000000000001001010100001", -- 4768 FREE #<CONS 0 4769>
 "00000000000000000001001010100010", -- 4769 FREE #<CONS 0 4770>
 "00000000000000000001001010100011", -- 4770 FREE #<CONS 0 4771>
 "00000000000000000001001010100100", -- 4771 FREE #<CONS 0 4772>
 "00000000000000000001001010100101", -- 4772 FREE #<CONS 0 4773>
 "00000000000000000001001010100110", -- 4773 FREE #<CONS 0 4774>
 "00000000000000000001001010100111", -- 4774 FREE #<CONS 0 4775>
 "00000000000000000001001010101000", -- 4775 FREE #<CONS 0 4776>
 "00000000000000000001001010101001", -- 4776 FREE #<CONS 0 4777>
 "00000000000000000001001010101010", -- 4777 FREE #<CONS 0 4778>
 "00000000000000000001001010101011", -- 4778 FREE #<CONS 0 4779>
 "00000000000000000001001010101100", -- 4779 FREE #<CONS 0 4780>
 "00000000000000000001001010101101", -- 4780 FREE #<CONS 0 4781>
 "00000000000000000001001010101110", -- 4781 FREE #<CONS 0 4782>
 "00000000000000000001001010101111", -- 4782 FREE #<CONS 0 4783>
 "00000000000000000001001010110000", -- 4783 FREE #<CONS 0 4784>
 "00000000000000000001001010110001", -- 4784 FREE #<CONS 0 4785>
 "00000000000000000001001010110010", -- 4785 FREE #<CONS 0 4786>
 "00000000000000000001001010110011", -- 4786 FREE #<CONS 0 4787>
 "00000000000000000001001010110100", -- 4787 FREE #<CONS 0 4788>
 "00000000000000000001001010110101", -- 4788 FREE #<CONS 0 4789>
 "00000000000000000001001010110110", -- 4789 FREE #<CONS 0 4790>
 "00000000000000000001001010110111", -- 4790 FREE #<CONS 0 4791>
 "00000000000000000001001010111000", -- 4791 FREE #<CONS 0 4792>
 "00000000000000000001001010111001", -- 4792 FREE #<CONS 0 4793>
 "00000000000000000001001010111010", -- 4793 FREE #<CONS 0 4794>
 "00000000000000000001001010111011", -- 4794 FREE #<CONS 0 4795>
 "00000000000000000001001010111100", -- 4795 FREE #<CONS 0 4796>
 "00000000000000000001001010111101", -- 4796 FREE #<CONS 0 4797>
 "00000000000000000001001010111110", -- 4797 FREE #<CONS 0 4798>
 "00000000000000000001001010111111", -- 4798 FREE #<CONS 0 4799>
 "00000000000000000001001011000000", -- 4799 FREE #<CONS 0 4800>
 "00000000000000000001001011000001", -- 4800 FREE #<CONS 0 4801>
 "00000000000000000001001011000010", -- 4801 FREE #<CONS 0 4802>
 "00000000000000000001001011000011", -- 4802 FREE #<CONS 0 4803>
 "00000000000000000001001011000100", -- 4803 FREE #<CONS 0 4804>
 "00000000000000000001001011000101", -- 4804 FREE #<CONS 0 4805>
 "00000000000000000001001011000110", -- 4805 FREE #<CONS 0 4806>
 "00000000000000000001001011000111", -- 4806 FREE #<CONS 0 4807>
 "00000000000000000001001011001000", -- 4807 FREE #<CONS 0 4808>
 "00000000000000000001001011001001", -- 4808 FREE #<CONS 0 4809>
 "00000000000000000001001011001010", -- 4809 FREE #<CONS 0 4810>
 "00000000000000000001001011001011", -- 4810 FREE #<CONS 0 4811>
 "00000000000000000001001011001100", -- 4811 FREE #<CONS 0 4812>
 "00000000000000000001001011001101", -- 4812 FREE #<CONS 0 4813>
 "00000000000000000001001011001110", -- 4813 FREE #<CONS 0 4814>
 "00000000000000000001001011001111", -- 4814 FREE #<CONS 0 4815>
 "00000000000000000001001011010000", -- 4815 FREE #<CONS 0 4816>
 "00000000000000000001001011010001", -- 4816 FREE #<CONS 0 4817>
 "00000000000000000001001011010010", -- 4817 FREE #<CONS 0 4818>
 "00000000000000000001001011010011", -- 4818 FREE #<CONS 0 4819>
 "00000000000000000001001011010100", -- 4819 FREE #<CONS 0 4820>
 "00000000000000000001001011010101", -- 4820 FREE #<CONS 0 4821>
 "00000000000000000001001011010110", -- 4821 FREE #<CONS 0 4822>
 "00000000000000000001001011010111", -- 4822 FREE #<CONS 0 4823>
 "00000000000000000001001011011000", -- 4823 FREE #<CONS 0 4824>
 "00000000000000000001001011011001", -- 4824 FREE #<CONS 0 4825>
 "00000000000000000001001011011010", -- 4825 FREE #<CONS 0 4826>
 "00000000000000000001001011011011", -- 4826 FREE #<CONS 0 4827>
 "00000000000000000001001011011100", -- 4827 FREE #<CONS 0 4828>
 "00000000000000000001001011011101", -- 4828 FREE #<CONS 0 4829>
 "00000000000000000001001011011110", -- 4829 FREE #<CONS 0 4830>
 "00000000000000000001001011011111", -- 4830 FREE #<CONS 0 4831>
 "00000000000000000001001011100000", -- 4831 FREE #<CONS 0 4832>
 "00000000000000000001001011100001", -- 4832 FREE #<CONS 0 4833>
 "00000000000000000001001011100010", -- 4833 FREE #<CONS 0 4834>
 "00000000000000000001001011100011", -- 4834 FREE #<CONS 0 4835>
 "00000000000000000001001011100100", -- 4835 FREE #<CONS 0 4836>
 "00000000000000000001001011100101", -- 4836 FREE #<CONS 0 4837>
 "00000000000000000001001011100110", -- 4837 FREE #<CONS 0 4838>
 "00000000000000000001001011100111", -- 4838 FREE #<CONS 0 4839>
 "00000000000000000001001011101000", -- 4839 FREE #<CONS 0 4840>
 "00000000000000000001001011101001", -- 4840 FREE #<CONS 0 4841>
 "00000000000000000001001011101010", -- 4841 FREE #<CONS 0 4842>
 "00000000000000000001001011101011", -- 4842 FREE #<CONS 0 4843>
 "00000000000000000001001011101100", -- 4843 FREE #<CONS 0 4844>
 "00000000000000000001001011101101", -- 4844 FREE #<CONS 0 4845>
 "00000000000000000001001011101110", -- 4845 FREE #<CONS 0 4846>
 "00000000000000000001001011101111", -- 4846 FREE #<CONS 0 4847>
 "00000000000000000001001011110000", -- 4847 FREE #<CONS 0 4848>
 "00000000000000000001001011110001", -- 4848 FREE #<CONS 0 4849>
 "00000000000000000001001011110010", -- 4849 FREE #<CONS 0 4850>
 "00000000000000000001001011110011", -- 4850 FREE #<CONS 0 4851>
 "00000000000000000001001011110100", -- 4851 FREE #<CONS 0 4852>
 "00000000000000000001001011110101", -- 4852 FREE #<CONS 0 4853>
 "00000000000000000001001011110110", -- 4853 FREE #<CONS 0 4854>
 "00000000000000000001001011110111", -- 4854 FREE #<CONS 0 4855>
 "00000000000000000001001011111000", -- 4855 FREE #<CONS 0 4856>
 "00000000000000000001001011111001", -- 4856 FREE #<CONS 0 4857>
 "00000000000000000001001011111010", -- 4857 FREE #<CONS 0 4858>
 "00000000000000000001001011111011", -- 4858 FREE #<CONS 0 4859>
 "00000000000000000001001011111100", -- 4859 FREE #<CONS 0 4860>
 "00000000000000000001001011111101", -- 4860 FREE #<CONS 0 4861>
 "00000000000000000001001011111110", -- 4861 FREE #<CONS 0 4862>
 "00000000000000000001001011111111", -- 4862 FREE #<CONS 0 4863>
 "00000000000000000001001100000000", -- 4863 FREE #<CONS 0 4864>
 "00000000000000000001001100000001", -- 4864 FREE #<CONS 0 4865>
 "00000000000000000001001100000010", -- 4865 FREE #<CONS 0 4866>
 "00000000000000000001001100000011", -- 4866 FREE #<CONS 0 4867>
 "00000000000000000001001100000100", -- 4867 FREE #<CONS 0 4868>
 "00000000000000000001001100000101", -- 4868 FREE #<CONS 0 4869>
 "00000000000000000001001100000110", -- 4869 FREE #<CONS 0 4870>
 "00000000000000000001001100000111", -- 4870 FREE #<CONS 0 4871>
 "00000000000000000001001100001000", -- 4871 FREE #<CONS 0 4872>
 "00000000000000000001001100001001", -- 4872 FREE #<CONS 0 4873>
 "00000000000000000001001100001010", -- 4873 FREE #<CONS 0 4874>
 "00000000000000000001001100001011", -- 4874 FREE #<CONS 0 4875>
 "00000000000000000001001100001100", -- 4875 FREE #<CONS 0 4876>
 "00000000000000000001001100001101", -- 4876 FREE #<CONS 0 4877>
 "00000000000000000001001100001110", -- 4877 FREE #<CONS 0 4878>
 "00000000000000000001001100001111", -- 4878 FREE #<CONS 0 4879>
 "00000000000000000001001100010000", -- 4879 FREE #<CONS 0 4880>
 "00000000000000000001001100010001", -- 4880 FREE #<CONS 0 4881>
 "00000000000000000001001100010010", -- 4881 FREE #<CONS 0 4882>
 "00000000000000000001001100010011", -- 4882 FREE #<CONS 0 4883>
 "00000000000000000001001100010100", -- 4883 FREE #<CONS 0 4884>
 "00000000000000000001001100010101", -- 4884 FREE #<CONS 0 4885>
 "00000000000000000001001100010110", -- 4885 FREE #<CONS 0 4886>
 "00000000000000000001001100010111", -- 4886 FREE #<CONS 0 4887>
 "00000000000000000001001100011000", -- 4887 FREE #<CONS 0 4888>
 "00000000000000000001001100011001", -- 4888 FREE #<CONS 0 4889>
 "00000000000000000001001100011010", -- 4889 FREE #<CONS 0 4890>
 "00000000000000000001001100011011", -- 4890 FREE #<CONS 0 4891>
 "00000000000000000001001100011100", -- 4891 FREE #<CONS 0 4892>
 "00000000000000000001001100011101", -- 4892 FREE #<CONS 0 4893>
 "00000000000000000001001100011110", -- 4893 FREE #<CONS 0 4894>
 "00000000000000000001001100011111", -- 4894 FREE #<CONS 0 4895>
 "00000000000000000001001100100000", -- 4895 FREE #<CONS 0 4896>
 "00000000000000000001001100100001", -- 4896 FREE #<CONS 0 4897>
 "00000000000000000001001100100010", -- 4897 FREE #<CONS 0 4898>
 "00000000000000000001001100100011", -- 4898 FREE #<CONS 0 4899>
 "00000000000000000001001100100100", -- 4899 FREE #<CONS 0 4900>
 "00000000000000000001001100100101", -- 4900 FREE #<CONS 0 4901>
 "00000000000000000001001100100110", -- 4901 FREE #<CONS 0 4902>
 "00000000000000000001001100100111", -- 4902 FREE #<CONS 0 4903>
 "00000000000000000001001100101000", -- 4903 FREE #<CONS 0 4904>
 "00000000000000000001001100101001", -- 4904 FREE #<CONS 0 4905>
 "00000000000000000001001100101010", -- 4905 FREE #<CONS 0 4906>
 "00000000000000000001001100101011", -- 4906 FREE #<CONS 0 4907>
 "00000000000000000001001100101100", -- 4907 FREE #<CONS 0 4908>
 "00000000000000000001001100101101", -- 4908 FREE #<CONS 0 4909>
 "00000000000000000001001100101110", -- 4909 FREE #<CONS 0 4910>
 "00000000000000000001001100101111", -- 4910 FREE #<CONS 0 4911>
 "00000000000000000001001100110000", -- 4911 FREE #<CONS 0 4912>
 "00000000000000000001001100110001", -- 4912 FREE #<CONS 0 4913>
 "00000000000000000001001100110010", -- 4913 FREE #<CONS 0 4914>
 "00000000000000000001001100110011", -- 4914 FREE #<CONS 0 4915>
 "00000000000000000001001100110100", -- 4915 FREE #<CONS 0 4916>
 "00000000000000000001001100110101", -- 4916 FREE #<CONS 0 4917>
 "00000000000000000001001100110110", -- 4917 FREE #<CONS 0 4918>
 "00000000000000000001001100110111", -- 4918 FREE #<CONS 0 4919>
 "00000000000000000001001100111000", -- 4919 FREE #<CONS 0 4920>
 "00000000000000000001001100111001", -- 4920 FREE #<CONS 0 4921>
 "00000000000000000001001100111010", -- 4921 FREE #<CONS 0 4922>
 "00000000000000000001001100111011", -- 4922 FREE #<CONS 0 4923>
 "00000000000000000001001100111100", -- 4923 FREE #<CONS 0 4924>
 "00000000000000000001001100111101", -- 4924 FREE #<CONS 0 4925>
 "00000000000000000001001100111110", -- 4925 FREE #<CONS 0 4926>
 "00000000000000000001001100111111", -- 4926 FREE #<CONS 0 4927>
 "00000000000000000001001101000000", -- 4927 FREE #<CONS 0 4928>
 "00000000000000000001001101000001", -- 4928 FREE #<CONS 0 4929>
 "00000000000000000001001101000010", -- 4929 FREE #<CONS 0 4930>
 "00000000000000000001001101000011", -- 4930 FREE #<CONS 0 4931>
 "00000000000000000001001101000100", -- 4931 FREE #<CONS 0 4932>
 "00000000000000000001001101000101", -- 4932 FREE #<CONS 0 4933>
 "00000000000000000001001101000110", -- 4933 FREE #<CONS 0 4934>
 "00000000000000000001001101000111", -- 4934 FREE #<CONS 0 4935>
 "00000000000000000001001101001000", -- 4935 FREE #<CONS 0 4936>
 "00000000000000000001001101001001", -- 4936 FREE #<CONS 0 4937>
 "00000000000000000001001101001010", -- 4937 FREE #<CONS 0 4938>
 "00000000000000000001001101001011", -- 4938 FREE #<CONS 0 4939>
 "00000000000000000001001101001100", -- 4939 FREE #<CONS 0 4940>
 "00000000000000000001001101001101", -- 4940 FREE #<CONS 0 4941>
 "00000000000000000001001101001110", -- 4941 FREE #<CONS 0 4942>
 "00000000000000000001001101001111", -- 4942 FREE #<CONS 0 4943>
 "00000000000000000001001101010000", -- 4943 FREE #<CONS 0 4944>
 "00000000000000000001001101010001", -- 4944 FREE #<CONS 0 4945>
 "00000000000000000001001101010010", -- 4945 FREE #<CONS 0 4946>
 "00000000000000000001001101010011", -- 4946 FREE #<CONS 0 4947>
 "00000000000000000001001101010100", -- 4947 FREE #<CONS 0 4948>
 "00000000000000000001001101010101", -- 4948 FREE #<CONS 0 4949>
 "00000000000000000001001101010110", -- 4949 FREE #<CONS 0 4950>
 "00000000000000000001001101010111", -- 4950 FREE #<CONS 0 4951>
 "00000000000000000001001101011000", -- 4951 FREE #<CONS 0 4952>
 "00000000000000000001001101011001", -- 4952 FREE #<CONS 0 4953>
 "00000000000000000001001101011010", -- 4953 FREE #<CONS 0 4954>
 "00000000000000000001001101011011", -- 4954 FREE #<CONS 0 4955>
 "00000000000000000001001101011100", -- 4955 FREE #<CONS 0 4956>
 "00000000000000000001001101011101", -- 4956 FREE #<CONS 0 4957>
 "00000000000000000001001101011110", -- 4957 FREE #<CONS 0 4958>
 "00000000000000000001001101011111", -- 4958 FREE #<CONS 0 4959>
 "00000000000000000001001101100000", -- 4959 FREE #<CONS 0 4960>
 "00000000000000000001001101100001", -- 4960 FREE #<CONS 0 4961>
 "00000000000000000001001101100010", -- 4961 FREE #<CONS 0 4962>
 "00000000000000000001001101100011", -- 4962 FREE #<CONS 0 4963>
 "00000000000000000001001101100100", -- 4963 FREE #<CONS 0 4964>
 "00000000000000000001001101100101", -- 4964 FREE #<CONS 0 4965>
 "00000000000000000001001101100110", -- 4965 FREE #<CONS 0 4966>
 "00000000000000000001001101100111", -- 4966 FREE #<CONS 0 4967>
 "00000000000000000001001101101000", -- 4967 FREE #<CONS 0 4968>
 "00000000000000000001001101101001", -- 4968 FREE #<CONS 0 4969>
 "00000000000000000001001101101010", -- 4969 FREE #<CONS 0 4970>
 "00000000000000000001001101101011", -- 4970 FREE #<CONS 0 4971>
 "00000000000000000001001101101100", -- 4971 FREE #<CONS 0 4972>
 "00000000000000000001001101101101", -- 4972 FREE #<CONS 0 4973>
 "00000000000000000001001101101110", -- 4973 FREE #<CONS 0 4974>
 "00000000000000000001001101101111", -- 4974 FREE #<CONS 0 4975>
 "00000000000000000001001101110000", -- 4975 FREE #<CONS 0 4976>
 "00000000000000000001001101110001", -- 4976 FREE #<CONS 0 4977>
 "00000000000000000001001101110010", -- 4977 FREE #<CONS 0 4978>
 "00000000000000000001001101110011", -- 4978 FREE #<CONS 0 4979>
 "00000000000000000001001101110100", -- 4979 FREE #<CONS 0 4980>
 "00000000000000000001001101110101", -- 4980 FREE #<CONS 0 4981>
 "00000000000000000001001101110110", -- 4981 FREE #<CONS 0 4982>
 "00000000000000000001001101110111", -- 4982 FREE #<CONS 0 4983>
 "00000000000000000001001101111000", -- 4983 FREE #<CONS 0 4984>
 "00000000000000000001001101111001", -- 4984 FREE #<CONS 0 4985>
 "00000000000000000001001101111010", -- 4985 FREE #<CONS 0 4986>
 "00000000000000000001001101111011", -- 4986 FREE #<CONS 0 4987>
 "00000000000000000001001101111100", -- 4987 FREE #<CONS 0 4988>
 "00000000000000000001001101111101", -- 4988 FREE #<CONS 0 4989>
 "00000000000000000001001101111110", -- 4989 FREE #<CONS 0 4990>
 "00000000000000000001001101111111", -- 4990 FREE #<CONS 0 4991>
 "00000000000000000001001110000000", -- 4991 FREE #<CONS 0 4992>
 "00000000000000000001001110000001", -- 4992 FREE #<CONS 0 4993>
 "00000000000000000001001110000010", -- 4993 FREE #<CONS 0 4994>
 "00000000000000000001001110000011", -- 4994 FREE #<CONS 0 4995>
 "00000000000000000001001110000100", -- 4995 FREE #<CONS 0 4996>
 "00000000000000000001001110000101", -- 4996 FREE #<CONS 0 4997>
 "00000000000000000001001110000110", -- 4997 FREE #<CONS 0 4998>
 "00000000000000000001001110000111", -- 4998 FREE #<CONS 0 4999>
 "00000000000000000001001110001000", -- 4999 FREE #<CONS 0 5000>
 "00000000000000000001001110001001", -- 5000 FREE #<CONS 0 5001>
 "00000000000000000001001110001010", -- 5001 FREE #<CONS 0 5002>
 "00000000000000000001001110001011", -- 5002 FREE #<CONS 0 5003>
 "00000000000000000001001110001100", -- 5003 FREE #<CONS 0 5004>
 "00000000000000000001001110001101", -- 5004 FREE #<CONS 0 5005>
 "00000000000000000001001110001110", -- 5005 FREE #<CONS 0 5006>
 "00000000000000000001001110001111", -- 5006 FREE #<CONS 0 5007>
 "00000000000000000001001110010000", -- 5007 FREE #<CONS 0 5008>
 "00000000000000000001001110010001", -- 5008 FREE #<CONS 0 5009>
 "00000000000000000001001110010010", -- 5009 FREE #<CONS 0 5010>
 "00000000000000000001001110010011", -- 5010 FREE #<CONS 0 5011>
 "00000000000000000001001110010100", -- 5011 FREE #<CONS 0 5012>
 "00000000000000000001001110010101", -- 5012 FREE #<CONS 0 5013>
 "00000000000000000001001110010110", -- 5013 FREE #<CONS 0 5014>
 "00000000000000000001001110010111", -- 5014 FREE #<CONS 0 5015>
 "00000000000000000001001110011000", -- 5015 FREE #<CONS 0 5016>
 "00000000000000000001001110011001", -- 5016 FREE #<CONS 0 5017>
 "00000000000000000001001110011010", -- 5017 FREE #<CONS 0 5018>
 "00000000000000000001001110011011", -- 5018 FREE #<CONS 0 5019>
 "00000000000000000001001110011100", -- 5019 FREE #<CONS 0 5020>
 "00000000000000000001001110011101", -- 5020 FREE #<CONS 0 5021>
 "00000000000000000001001110011110", -- 5021 FREE #<CONS 0 5022>
 "00000000000000000001001110011111", -- 5022 FREE #<CONS 0 5023>
 "00000000000000000001001110100000", -- 5023 FREE #<CONS 0 5024>
 "00000000000000000001001110100001", -- 5024 FREE #<CONS 0 5025>
 "00000000000000000001001110100010", -- 5025 FREE #<CONS 0 5026>
 "00000000000000000001001110100011", -- 5026 FREE #<CONS 0 5027>
 "00000000000000000001001110100100", -- 5027 FREE #<CONS 0 5028>
 "00000000000000000001001110100101", -- 5028 FREE #<CONS 0 5029>
 "00000000000000000001001110100110", -- 5029 FREE #<CONS 0 5030>
 "00000000000000000001001110100111", -- 5030 FREE #<CONS 0 5031>
 "00000000000000000001001110101000", -- 5031 FREE #<CONS 0 5032>
 "00000000000000000001001110101001", -- 5032 FREE #<CONS 0 5033>
 "00000000000000000001001110101010", -- 5033 FREE #<CONS 0 5034>
 "00000000000000000001001110101011", -- 5034 FREE #<CONS 0 5035>
 "00000000000000000001001110101100", -- 5035 FREE #<CONS 0 5036>
 "00000000000000000001001110101101", -- 5036 FREE #<CONS 0 5037>
 "00000000000000000001001110101110", -- 5037 FREE #<CONS 0 5038>
 "00000000000000000001001110101111", -- 5038 FREE #<CONS 0 5039>
 "00000000000000000001001110110000", -- 5039 FREE #<CONS 0 5040>
 "00000000000000000001001110110001", -- 5040 FREE #<CONS 0 5041>
 "00000000000000000001001110110010", -- 5041 FREE #<CONS 0 5042>
 "00000000000000000001001110110011", -- 5042 FREE #<CONS 0 5043>
 "00000000000000000001001110110100", -- 5043 FREE #<CONS 0 5044>
 "00000000000000000001001110110101", -- 5044 FREE #<CONS 0 5045>
 "00000000000000000001001110110110", -- 5045 FREE #<CONS 0 5046>
 "00000000000000000001001110110111", -- 5046 FREE #<CONS 0 5047>
 "00000000000000000001001110111000", -- 5047 FREE #<CONS 0 5048>
 "00000000000000000001001110111001", -- 5048 FREE #<CONS 0 5049>
 "00000000000000000001001110111010", -- 5049 FREE #<CONS 0 5050>
 "00000000000000000001001110111011", -- 5050 FREE #<CONS 0 5051>
 "00000000000000000001001110111100", -- 5051 FREE #<CONS 0 5052>
 "00000000000000000001001110111101", -- 5052 FREE #<CONS 0 5053>
 "00000000000000000001001110111110", -- 5053 FREE #<CONS 0 5054>
 "00000000000000000001001110111111", -- 5054 FREE #<CONS 0 5055>
 "00000000000000000001001111000000", -- 5055 FREE #<CONS 0 5056>
 "00000000000000000001001111000001", -- 5056 FREE #<CONS 0 5057>
 "00000000000000000001001111000010", -- 5057 FREE #<CONS 0 5058>
 "00000000000000000001001111000011", -- 5058 FREE #<CONS 0 5059>
 "00000000000000000001001111000100", -- 5059 FREE #<CONS 0 5060>
 "00000000000000000001001111000101", -- 5060 FREE #<CONS 0 5061>
 "00000000000000000001001111000110", -- 5061 FREE #<CONS 0 5062>
 "00000000000000000001001111000111", -- 5062 FREE #<CONS 0 5063>
 "00000000000000000001001111001000", -- 5063 FREE #<CONS 0 5064>
 "00000000000000000001001111001001", -- 5064 FREE #<CONS 0 5065>
 "00000000000000000001001111001010", -- 5065 FREE #<CONS 0 5066>
 "00000000000000000001001111001011", -- 5066 FREE #<CONS 0 5067>
 "00000000000000000001001111001100", -- 5067 FREE #<CONS 0 5068>
 "00000000000000000001001111001101", -- 5068 FREE #<CONS 0 5069>
 "00000000000000000001001111001110", -- 5069 FREE #<CONS 0 5070>
 "00000000000000000001001111001111", -- 5070 FREE #<CONS 0 5071>
 "00000000000000000001001111010000", -- 5071 FREE #<CONS 0 5072>
 "00000000000000000001001111010001", -- 5072 FREE #<CONS 0 5073>
 "00000000000000000001001111010010", -- 5073 FREE #<CONS 0 5074>
 "00000000000000000001001111010011", -- 5074 FREE #<CONS 0 5075>
 "00000000000000000001001111010100", -- 5075 FREE #<CONS 0 5076>
 "00000000000000000001001111010101", -- 5076 FREE #<CONS 0 5077>
 "00000000000000000001001111010110", -- 5077 FREE #<CONS 0 5078>
 "00000000000000000001001111010111", -- 5078 FREE #<CONS 0 5079>
 "00000000000000000001001111011000", -- 5079 FREE #<CONS 0 5080>
 "00000000000000000001001111011001", -- 5080 FREE #<CONS 0 5081>
 "00000000000000000001001111011010", -- 5081 FREE #<CONS 0 5082>
 "00000000000000000001001111011011", -- 5082 FREE #<CONS 0 5083>
 "00000000000000000001001111011100", -- 5083 FREE #<CONS 0 5084>
 "00000000000000000001001111011101", -- 5084 FREE #<CONS 0 5085>
 "00000000000000000001001111011110", -- 5085 FREE #<CONS 0 5086>
 "00000000000000000001001111011111", -- 5086 FREE #<CONS 0 5087>
 "00000000000000000001001111100000", -- 5087 FREE #<CONS 0 5088>
 "00000000000000000001001111100001", -- 5088 FREE #<CONS 0 5089>
 "00000000000000000001001111100010", -- 5089 FREE #<CONS 0 5090>
 "00000000000000000001001111100011", -- 5090 FREE #<CONS 0 5091>
 "00000000000000000001001111100100", -- 5091 FREE #<CONS 0 5092>
 "00000000000000000001001111100101", -- 5092 FREE #<CONS 0 5093>
 "00000000000000000001001111100110", -- 5093 FREE #<CONS 0 5094>
 "00000000000000000001001111100111", -- 5094 FREE #<CONS 0 5095>
 "00000000000000000001001111101000", -- 5095 FREE #<CONS 0 5096>
 "00000000000000000001001111101001", -- 5096 FREE #<CONS 0 5097>
 "00000000000000000001001111101010", -- 5097 FREE #<CONS 0 5098>
 "00000000000000000001001111101011", -- 5098 FREE #<CONS 0 5099>
 "00000000000000000001001111101100", -- 5099 FREE #<CONS 0 5100>
 "00000000000000000001001111101101", -- 5100 FREE #<CONS 0 5101>
 "00000000000000000001001111101110", -- 5101 FREE #<CONS 0 5102>
 "00000000000000000001001111101111", -- 5102 FREE #<CONS 0 5103>
 "00000000000000000001001111110000", -- 5103 FREE #<CONS 0 5104>
 "00000000000000000001001111110001", -- 5104 FREE #<CONS 0 5105>
 "00000000000000000001001111110010", -- 5105 FREE #<CONS 0 5106>
 "00000000000000000001001111110011", -- 5106 FREE #<CONS 0 5107>
 "00000000000000000001001111110100", -- 5107 FREE #<CONS 0 5108>
 "00000000000000000001001111110101", -- 5108 FREE #<CONS 0 5109>
 "00000000000000000001001111110110", -- 5109 FREE #<CONS 0 5110>
 "00000000000000000001001111110111", -- 5110 FREE #<CONS 0 5111>
 "00000000000000000001001111111000", -- 5111 FREE #<CONS 0 5112>
 "00000000000000000001001111111001", -- 5112 FREE #<CONS 0 5113>
 "00000000000000000001001111111010", -- 5113 FREE #<CONS 0 5114>
 "00000000000000000001001111111011", -- 5114 FREE #<CONS 0 5115>
 "00000000000000000001001111111100", -- 5115 FREE #<CONS 0 5116>
 "00000000000000000001001111111101", -- 5116 FREE #<CONS 0 5117>
 "00000000000000000001001111111110", -- 5117 FREE #<CONS 0 5118>
 "00000000000000000001001111111111", -- 5118 FREE #<CONS 0 5119>
 "00000000000000000001010000000000", -- 5119 FREE #<CONS 0 5120>
 "00000000000000000001010000000001", -- 5120 FREE #<CONS 0 5121>
 "00000000000000000001010000000010", -- 5121 FREE #<CONS 0 5122>
 "00000000000000000001010000000011", -- 5122 FREE #<CONS 0 5123>
 "00000000000000000001010000000100", -- 5123 FREE #<CONS 0 5124>
 "00000000000000000001010000000101", -- 5124 FREE #<CONS 0 5125>
 "00000000000000000001010000000110", -- 5125 FREE #<CONS 0 5126>
 "00000000000000000001010000000111", -- 5126 FREE #<CONS 0 5127>
 "00000000000000000001010000001000", -- 5127 FREE #<CONS 0 5128>
 "00000000000000000001010000001001", -- 5128 FREE #<CONS 0 5129>
 "00000000000000000001010000001010", -- 5129 FREE #<CONS 0 5130>
 "00000000000000000001010000001011", -- 5130 FREE #<CONS 0 5131>
 "00000000000000000001010000001100", -- 5131 FREE #<CONS 0 5132>
 "00000000000000000001010000001101", -- 5132 FREE #<CONS 0 5133>
 "00000000000000000001010000001110", -- 5133 FREE #<CONS 0 5134>
 "00000000000000000001010000001111", -- 5134 FREE #<CONS 0 5135>
 "00000000000000000001010000010000", -- 5135 FREE #<CONS 0 5136>
 "00000000000000000001010000010001", -- 5136 FREE #<CONS 0 5137>
 "00000000000000000001010000010010", -- 5137 FREE #<CONS 0 5138>
 "00000000000000000001010000010011", -- 5138 FREE #<CONS 0 5139>
 "00000000000000000001010000010100", -- 5139 FREE #<CONS 0 5140>
 "00000000000000000001010000010101", -- 5140 FREE #<CONS 0 5141>
 "00000000000000000001010000010110", -- 5141 FREE #<CONS 0 5142>
 "00000000000000000001010000010111", -- 5142 FREE #<CONS 0 5143>
 "00000000000000000001010000011000", -- 5143 FREE #<CONS 0 5144>
 "00000000000000000001010000011001", -- 5144 FREE #<CONS 0 5145>
 "00000000000000000001010000011010", -- 5145 FREE #<CONS 0 5146>
 "00000000000000000001010000011011", -- 5146 FREE #<CONS 0 5147>
 "00000000000000000001010000011100", -- 5147 FREE #<CONS 0 5148>
 "00000000000000000001010000011101", -- 5148 FREE #<CONS 0 5149>
 "00000000000000000001010000011110", -- 5149 FREE #<CONS 0 5150>
 "00000000000000000001010000011111", -- 5150 FREE #<CONS 0 5151>
 "00000000000000000001010000100000", -- 5151 FREE #<CONS 0 5152>
 "00000000000000000001010000100001", -- 5152 FREE #<CONS 0 5153>
 "00000000000000000001010000100010", -- 5153 FREE #<CONS 0 5154>
 "00000000000000000001010000100011", -- 5154 FREE #<CONS 0 5155>
 "00000000000000000001010000100100", -- 5155 FREE #<CONS 0 5156>
 "00000000000000000001010000100101", -- 5156 FREE #<CONS 0 5157>
 "00000000000000000001010000100110", -- 5157 FREE #<CONS 0 5158>
 "00000000000000000001010000100111", -- 5158 FREE #<CONS 0 5159>
 "00000000000000000001010000101000", -- 5159 FREE #<CONS 0 5160>
 "00000000000000000001010000101001", -- 5160 FREE #<CONS 0 5161>
 "00000000000000000001010000101010", -- 5161 FREE #<CONS 0 5162>
 "00000000000000000001010000101011", -- 5162 FREE #<CONS 0 5163>
 "00000000000000000001010000101100", -- 5163 FREE #<CONS 0 5164>
 "00000000000000000001010000101101", -- 5164 FREE #<CONS 0 5165>
 "00000000000000000001010000101110", -- 5165 FREE #<CONS 0 5166>
 "00000000000000000001010000101111", -- 5166 FREE #<CONS 0 5167>
 "00000000000000000001010000110000", -- 5167 FREE #<CONS 0 5168>
 "00000000000000000001010000110001", -- 5168 FREE #<CONS 0 5169>
 "00000000000000000001010000110010", -- 5169 FREE #<CONS 0 5170>
 "00000000000000000001010000110011", -- 5170 FREE #<CONS 0 5171>
 "00000000000000000001010000110100", -- 5171 FREE #<CONS 0 5172>
 "00000000000000000001010000110101", -- 5172 FREE #<CONS 0 5173>
 "00000000000000000001010000110110", -- 5173 FREE #<CONS 0 5174>
 "00000000000000000001010000110111", -- 5174 FREE #<CONS 0 5175>
 "00000000000000000001010000111000", -- 5175 FREE #<CONS 0 5176>
 "00000000000000000001010000111001", -- 5176 FREE #<CONS 0 5177>
 "00000000000000000001010000111010", -- 5177 FREE #<CONS 0 5178>
 "00000000000000000001010000111011", -- 5178 FREE #<CONS 0 5179>
 "00000000000000000001010000111100", -- 5179 FREE #<CONS 0 5180>
 "00000000000000000001010000111101", -- 5180 FREE #<CONS 0 5181>
 "00000000000000000001010000111110", -- 5181 FREE #<CONS 0 5182>
 "00000000000000000001010000111111", -- 5182 FREE #<CONS 0 5183>
 "00000000000000000001010001000000", -- 5183 FREE #<CONS 0 5184>
 "00000000000000000001010001000001", -- 5184 FREE #<CONS 0 5185>
 "00000000000000000001010001000010", -- 5185 FREE #<CONS 0 5186>
 "00000000000000000001010001000011", -- 5186 FREE #<CONS 0 5187>
 "00000000000000000001010001000100", -- 5187 FREE #<CONS 0 5188>
 "00000000000000000001010001000101", -- 5188 FREE #<CONS 0 5189>
 "00000000000000000001010001000110", -- 5189 FREE #<CONS 0 5190>
 "00000000000000000001010001000111", -- 5190 FREE #<CONS 0 5191>
 "00000000000000000001010001001000", -- 5191 FREE #<CONS 0 5192>
 "00000000000000000001010001001001", -- 5192 FREE #<CONS 0 5193>
 "00000000000000000001010001001010", -- 5193 FREE #<CONS 0 5194>
 "00000000000000000001010001001011", -- 5194 FREE #<CONS 0 5195>
 "00000000000000000001010001001100", -- 5195 FREE #<CONS 0 5196>
 "00000000000000000001010001001101", -- 5196 FREE #<CONS 0 5197>
 "00000000000000000001010001001110", -- 5197 FREE #<CONS 0 5198>
 "00000000000000000001010001001111", -- 5198 FREE #<CONS 0 5199>
 "00000000000000000001010001010000", -- 5199 FREE #<CONS 0 5200>
 "00000000000000000001010001010001", -- 5200 FREE #<CONS 0 5201>
 "00000000000000000001010001010010", -- 5201 FREE #<CONS 0 5202>
 "00000000000000000001010001010011", -- 5202 FREE #<CONS 0 5203>
 "00000000000000000001010001010100", -- 5203 FREE #<CONS 0 5204>
 "00000000000000000001010001010101", -- 5204 FREE #<CONS 0 5205>
 "00000000000000000001010001010110", -- 5205 FREE #<CONS 0 5206>
 "00000000000000000001010001010111", -- 5206 FREE #<CONS 0 5207>
 "00000000000000000001010001011000", -- 5207 FREE #<CONS 0 5208>
 "00000000000000000001010001011001", -- 5208 FREE #<CONS 0 5209>
 "00000000000000000001010001011010", -- 5209 FREE #<CONS 0 5210>
 "00000000000000000001010001011011", -- 5210 FREE #<CONS 0 5211>
 "00000000000000000001010001011100", -- 5211 FREE #<CONS 0 5212>
 "00000000000000000001010001011101", -- 5212 FREE #<CONS 0 5213>
 "00000000000000000001010001011110", -- 5213 FREE #<CONS 0 5214>
 "00000000000000000001010001011111", -- 5214 FREE #<CONS 0 5215>
 "00000000000000000001010001100000", -- 5215 FREE #<CONS 0 5216>
 "00000000000000000001010001100001", -- 5216 FREE #<CONS 0 5217>
 "00000000000000000001010001100010", -- 5217 FREE #<CONS 0 5218>
 "00000000000000000001010001100011", -- 5218 FREE #<CONS 0 5219>
 "00000000000000000001010001100100", -- 5219 FREE #<CONS 0 5220>
 "00000000000000000001010001100101", -- 5220 FREE #<CONS 0 5221>
 "00000000000000000001010001100110", -- 5221 FREE #<CONS 0 5222>
 "00000000000000000001010001100111", -- 5222 FREE #<CONS 0 5223>
 "00000000000000000001010001101000", -- 5223 FREE #<CONS 0 5224>
 "00000000000000000001010001101001", -- 5224 FREE #<CONS 0 5225>
 "00000000000000000001010001101010", -- 5225 FREE #<CONS 0 5226>
 "00000000000000000001010001101011", -- 5226 FREE #<CONS 0 5227>
 "00000000000000000001010001101100", -- 5227 FREE #<CONS 0 5228>
 "00000000000000000001010001101101", -- 5228 FREE #<CONS 0 5229>
 "00000000000000000001010001101110", -- 5229 FREE #<CONS 0 5230>
 "00000000000000000001010001101111", -- 5230 FREE #<CONS 0 5231>
 "00000000000000000001010001110000", -- 5231 FREE #<CONS 0 5232>
 "00000000000000000001010001110001", -- 5232 FREE #<CONS 0 5233>
 "00000000000000000001010001110010", -- 5233 FREE #<CONS 0 5234>
 "00000000000000000001010001110011", -- 5234 FREE #<CONS 0 5235>
 "00000000000000000001010001110100", -- 5235 FREE #<CONS 0 5236>
 "00000000000000000001010001110101", -- 5236 FREE #<CONS 0 5237>
 "00000000000000000001010001110110", -- 5237 FREE #<CONS 0 5238>
 "00000000000000000001010001110111", -- 5238 FREE #<CONS 0 5239>
 "00000000000000000001010001111000", -- 5239 FREE #<CONS 0 5240>
 "00000000000000000001010001111001", -- 5240 FREE #<CONS 0 5241>
 "00000000000000000001010001111010", -- 5241 FREE #<CONS 0 5242>
 "00000000000000000001010001111011", -- 5242 FREE #<CONS 0 5243>
 "00000000000000000001010001111100", -- 5243 FREE #<CONS 0 5244>
 "00000000000000000001010001111101", -- 5244 FREE #<CONS 0 5245>
 "00000000000000000001010001111110", -- 5245 FREE #<CONS 0 5246>
 "00000000000000000001010001111111", -- 5246 FREE #<CONS 0 5247>
 "00000000000000000001010010000000", -- 5247 FREE #<CONS 0 5248>
 "00000000000000000001010010000001", -- 5248 FREE #<CONS 0 5249>
 "00000000000000000001010010000010", -- 5249 FREE #<CONS 0 5250>
 "00000000000000000001010010000011", -- 5250 FREE #<CONS 0 5251>
 "00000000000000000001010010000100", -- 5251 FREE #<CONS 0 5252>
 "00000000000000000001010010000101", -- 5252 FREE #<CONS 0 5253>
 "00000000000000000001010010000110", -- 5253 FREE #<CONS 0 5254>
 "00000000000000000001010010000111", -- 5254 FREE #<CONS 0 5255>
 "00000000000000000001010010001000", -- 5255 FREE #<CONS 0 5256>
 "00000000000000000001010010001001", -- 5256 FREE #<CONS 0 5257>
 "00000000000000000001010010001010", -- 5257 FREE #<CONS 0 5258>
 "00000000000000000001010010001011", -- 5258 FREE #<CONS 0 5259>
 "00000000000000000001010010001100", -- 5259 FREE #<CONS 0 5260>
 "00000000000000000001010010001101", -- 5260 FREE #<CONS 0 5261>
 "00000000000000000001010010001110", -- 5261 FREE #<CONS 0 5262>
 "00000000000000000001010010001111", -- 5262 FREE #<CONS 0 5263>
 "00000000000000000001010010010000", -- 5263 FREE #<CONS 0 5264>
 "00000000000000000001010010010001", -- 5264 FREE #<CONS 0 5265>
 "00000000000000000001010010010010", -- 5265 FREE #<CONS 0 5266>
 "00000000000000000001010010010011", -- 5266 FREE #<CONS 0 5267>
 "00000000000000000001010010010100", -- 5267 FREE #<CONS 0 5268>
 "00000000000000000001010010010101", -- 5268 FREE #<CONS 0 5269>
 "00000000000000000001010010010110", -- 5269 FREE #<CONS 0 5270>
 "00000000000000000001010010010111", -- 5270 FREE #<CONS 0 5271>
 "00000000000000000001010010011000", -- 5271 FREE #<CONS 0 5272>
 "00000000000000000001010010011001", -- 5272 FREE #<CONS 0 5273>
 "00000000000000000001010010011010", -- 5273 FREE #<CONS 0 5274>
 "00000000000000000001010010011011", -- 5274 FREE #<CONS 0 5275>
 "00000000000000000001010010011100", -- 5275 FREE #<CONS 0 5276>
 "00000000000000000001010010011101", -- 5276 FREE #<CONS 0 5277>
 "00000000000000000001010010011110", -- 5277 FREE #<CONS 0 5278>
 "00000000000000000001010010011111", -- 5278 FREE #<CONS 0 5279>
 "00000000000000000001010010100000", -- 5279 FREE #<CONS 0 5280>
 "00000000000000000001010010100001", -- 5280 FREE #<CONS 0 5281>
 "00000000000000000001010010100010", -- 5281 FREE #<CONS 0 5282>
 "00000000000000000001010010100011", -- 5282 FREE #<CONS 0 5283>
 "00000000000000000001010010100100", -- 5283 FREE #<CONS 0 5284>
 "00000000000000000001010010100101", -- 5284 FREE #<CONS 0 5285>
 "00000000000000000001010010100110", -- 5285 FREE #<CONS 0 5286>
 "00000000000000000001010010100111", -- 5286 FREE #<CONS 0 5287>
 "00000000000000000001010010101000", -- 5287 FREE #<CONS 0 5288>
 "00000000000000000001010010101001", -- 5288 FREE #<CONS 0 5289>
 "00000000000000000001010010101010", -- 5289 FREE #<CONS 0 5290>
 "00000000000000000001010010101011", -- 5290 FREE #<CONS 0 5291>
 "00000000000000000001010010101100", -- 5291 FREE #<CONS 0 5292>
 "00000000000000000001010010101101", -- 5292 FREE #<CONS 0 5293>
 "00000000000000000001010010101110", -- 5293 FREE #<CONS 0 5294>
 "00000000000000000001010010101111", -- 5294 FREE #<CONS 0 5295>
 "00000000000000000001010010110000", -- 5295 FREE #<CONS 0 5296>
 "00000000000000000001010010110001", -- 5296 FREE #<CONS 0 5297>
 "00000000000000000001010010110010", -- 5297 FREE #<CONS 0 5298>
 "00000000000000000001010010110011", -- 5298 FREE #<CONS 0 5299>
 "00000000000000000001010010110100", -- 5299 FREE #<CONS 0 5300>
 "00000000000000000001010010110101", -- 5300 FREE #<CONS 0 5301>
 "00000000000000000001010010110110", -- 5301 FREE #<CONS 0 5302>
 "00000000000000000001010010110111", -- 5302 FREE #<CONS 0 5303>
 "00000000000000000001010010111000", -- 5303 FREE #<CONS 0 5304>
 "00000000000000000001010010111001", -- 5304 FREE #<CONS 0 5305>
 "00000000000000000001010010111010", -- 5305 FREE #<CONS 0 5306>
 "00000000000000000001010010111011", -- 5306 FREE #<CONS 0 5307>
 "00000000000000000001010010111100", -- 5307 FREE #<CONS 0 5308>
 "00000000000000000001010010111101", -- 5308 FREE #<CONS 0 5309>
 "00000000000000000001010010111110", -- 5309 FREE #<CONS 0 5310>
 "00000000000000000001010010111111", -- 5310 FREE #<CONS 0 5311>
 "00000000000000000001010011000000", -- 5311 FREE #<CONS 0 5312>
 "00000000000000000001010011000001", -- 5312 FREE #<CONS 0 5313>
 "00000000000000000001010011000010", -- 5313 FREE #<CONS 0 5314>
 "00000000000000000001010011000011", -- 5314 FREE #<CONS 0 5315>
 "00000000000000000001010011000100", -- 5315 FREE #<CONS 0 5316>
 "00000000000000000001010011000101", -- 5316 FREE #<CONS 0 5317>
 "00000000000000000001010011000110", -- 5317 FREE #<CONS 0 5318>
 "00000000000000000001010011000111", -- 5318 FREE #<CONS 0 5319>
 "00000000000000000001010011001000", -- 5319 FREE #<CONS 0 5320>
 "00000000000000000001010011001001", -- 5320 FREE #<CONS 0 5321>
 "00000000000000000001010011001010", -- 5321 FREE #<CONS 0 5322>
 "00000000000000000001010011001011", -- 5322 FREE #<CONS 0 5323>
 "00000000000000000001010011001100", -- 5323 FREE #<CONS 0 5324>
 "00000000000000000001010011001101", -- 5324 FREE #<CONS 0 5325>
 "00000000000000000001010011001110", -- 5325 FREE #<CONS 0 5326>
 "00000000000000000001010011001111", -- 5326 FREE #<CONS 0 5327>
 "00000000000000000001010011010000", -- 5327 FREE #<CONS 0 5328>
 "00000000000000000001010011010001", -- 5328 FREE #<CONS 0 5329>
 "00000000000000000001010011010010", -- 5329 FREE #<CONS 0 5330>
 "00000000000000000001010011010011", -- 5330 FREE #<CONS 0 5331>
 "00000000000000000001010011010100", -- 5331 FREE #<CONS 0 5332>
 "00000000000000000001010011010101", -- 5332 FREE #<CONS 0 5333>
 "00000000000000000001010011010110", -- 5333 FREE #<CONS 0 5334>
 "00000000000000000001010011010111", -- 5334 FREE #<CONS 0 5335>
 "00000000000000000001010011011000", -- 5335 FREE #<CONS 0 5336>
 "00000000000000000001010011011001", -- 5336 FREE #<CONS 0 5337>
 "00000000000000000001010011011010", -- 5337 FREE #<CONS 0 5338>
 "00000000000000000001010011011011", -- 5338 FREE #<CONS 0 5339>
 "00000000000000000001010011011100", -- 5339 FREE #<CONS 0 5340>
 "00000000000000000001010011011101", -- 5340 FREE #<CONS 0 5341>
 "00000000000000000001010011011110", -- 5341 FREE #<CONS 0 5342>
 "00000000000000000001010011011111", -- 5342 FREE #<CONS 0 5343>
 "00000000000000000001010011100000", -- 5343 FREE #<CONS 0 5344>
 "00000000000000000001010011100001", -- 5344 FREE #<CONS 0 5345>
 "00000000000000000001010011100010", -- 5345 FREE #<CONS 0 5346>
 "00000000000000000001010011100011", -- 5346 FREE #<CONS 0 5347>
 "00000000000000000001010011100100", -- 5347 FREE #<CONS 0 5348>
 "00000000000000000001010011100101", -- 5348 FREE #<CONS 0 5349>
 "00000000000000000001010011100110", -- 5349 FREE #<CONS 0 5350>
 "00000000000000000001010011100111", -- 5350 FREE #<CONS 0 5351>
 "00000000000000000001010011101000", -- 5351 FREE #<CONS 0 5352>
 "00000000000000000001010011101001", -- 5352 FREE #<CONS 0 5353>
 "00000000000000000001010011101010", -- 5353 FREE #<CONS 0 5354>
 "00000000000000000001010011101011", -- 5354 FREE #<CONS 0 5355>
 "00000000000000000001010011101100", -- 5355 FREE #<CONS 0 5356>
 "00000000000000000001010011101101", -- 5356 FREE #<CONS 0 5357>
 "00000000000000000001010011101110", -- 5357 FREE #<CONS 0 5358>
 "00000000000000000001010011101111", -- 5358 FREE #<CONS 0 5359>
 "00000000000000000001010011110000", -- 5359 FREE #<CONS 0 5360>
 "00000000000000000001010011110001", -- 5360 FREE #<CONS 0 5361>
 "00000000000000000001010011110010", -- 5361 FREE #<CONS 0 5362>
 "00000000000000000001010011110011", -- 5362 FREE #<CONS 0 5363>
 "00000000000000000001010011110100", -- 5363 FREE #<CONS 0 5364>
 "00000000000000000001010011110101", -- 5364 FREE #<CONS 0 5365>
 "00000000000000000001010011110110", -- 5365 FREE #<CONS 0 5366>
 "00000000000000000001010011110111", -- 5366 FREE #<CONS 0 5367>
 "00000000000000000001010011111000", -- 5367 FREE #<CONS 0 5368>
 "00000000000000000001010011111001", -- 5368 FREE #<CONS 0 5369>
 "00000000000000000001010011111010", -- 5369 FREE #<CONS 0 5370>
 "00000000000000000001010011111011", -- 5370 FREE #<CONS 0 5371>
 "00000000000000000001010011111100", -- 5371 FREE #<CONS 0 5372>
 "00000000000000000001010011111101", -- 5372 FREE #<CONS 0 5373>
 "00000000000000000001010011111110", -- 5373 FREE #<CONS 0 5374>
 "00000000000000000001010011111111", -- 5374 FREE #<CONS 0 5375>
 "00000000000000000001010100000000", -- 5375 FREE #<CONS 0 5376>
 "00000000000000000001010100000001", -- 5376 FREE #<CONS 0 5377>
 "00000000000000000001010100000010", -- 5377 FREE #<CONS 0 5378>
 "00000000000000000001010100000011", -- 5378 FREE #<CONS 0 5379>
 "00000000000000000001010100000100", -- 5379 FREE #<CONS 0 5380>
 "00000000000000000001010100000101", -- 5380 FREE #<CONS 0 5381>
 "00000000000000000001010100000110", -- 5381 FREE #<CONS 0 5382>
 "00000000000000000001010100000111", -- 5382 FREE #<CONS 0 5383>
 "00000000000000000001010100001000", -- 5383 FREE #<CONS 0 5384>
 "00000000000000000001010100001001", -- 5384 FREE #<CONS 0 5385>
 "00000000000000000001010100001010", -- 5385 FREE #<CONS 0 5386>
 "00000000000000000001010100001011", -- 5386 FREE #<CONS 0 5387>
 "00000000000000000001010100001100", -- 5387 FREE #<CONS 0 5388>
 "00000000000000000001010100001101", -- 5388 FREE #<CONS 0 5389>
 "00000000000000000001010100001110", -- 5389 FREE #<CONS 0 5390>
 "00000000000000000001010100001111", -- 5390 FREE #<CONS 0 5391>
 "00000000000000000001010100010000", -- 5391 FREE #<CONS 0 5392>
 "00000000000000000001010100010001", -- 5392 FREE #<CONS 0 5393>
 "00000000000000000001010100010010", -- 5393 FREE #<CONS 0 5394>
 "00000000000000000001010100010011", -- 5394 FREE #<CONS 0 5395>
 "00000000000000000001010100010100", -- 5395 FREE #<CONS 0 5396>
 "00000000000000000001010100010101", -- 5396 FREE #<CONS 0 5397>
 "00000000000000000001010100010110", -- 5397 FREE #<CONS 0 5398>
 "00000000000000000001010100010111", -- 5398 FREE #<CONS 0 5399>
 "00000000000000000001010100011000", -- 5399 FREE #<CONS 0 5400>
 "00000000000000000001010100011001", -- 5400 FREE #<CONS 0 5401>
 "00000000000000000001010100011010", -- 5401 FREE #<CONS 0 5402>
 "00000000000000000001010100011011", -- 5402 FREE #<CONS 0 5403>
 "00000000000000000001010100011100", -- 5403 FREE #<CONS 0 5404>
 "00000000000000000001010100011101", -- 5404 FREE #<CONS 0 5405>
 "00000000000000000001010100011110", -- 5405 FREE #<CONS 0 5406>
 "00000000000000000001010100011111", -- 5406 FREE #<CONS 0 5407>
 "00000000000000000001010100100000", -- 5407 FREE #<CONS 0 5408>
 "00000000000000000001010100100001", -- 5408 FREE #<CONS 0 5409>
 "00000000000000000001010100100010", -- 5409 FREE #<CONS 0 5410>
 "00000000000000000001010100100011", -- 5410 FREE #<CONS 0 5411>
 "00000000000000000001010100100100", -- 5411 FREE #<CONS 0 5412>
 "00000000000000000001010100100101", -- 5412 FREE #<CONS 0 5413>
 "00000000000000000001010100100110", -- 5413 FREE #<CONS 0 5414>
 "00000000000000000001010100100111", -- 5414 FREE #<CONS 0 5415>
 "00000000000000000001010100101000", -- 5415 FREE #<CONS 0 5416>
 "00000000000000000001010100101001", -- 5416 FREE #<CONS 0 5417>
 "00000000000000000001010100101010", -- 5417 FREE #<CONS 0 5418>
 "00000000000000000001010100101011", -- 5418 FREE #<CONS 0 5419>
 "00000000000000000001010100101100", -- 5419 FREE #<CONS 0 5420>
 "00000000000000000001010100101101", -- 5420 FREE #<CONS 0 5421>
 "00000000000000000001010100101110", -- 5421 FREE #<CONS 0 5422>
 "00000000000000000001010100101111", -- 5422 FREE #<CONS 0 5423>
 "00000000000000000001010100110000", -- 5423 FREE #<CONS 0 5424>
 "00000000000000000001010100110001", -- 5424 FREE #<CONS 0 5425>
 "00000000000000000001010100110010", -- 5425 FREE #<CONS 0 5426>
 "00000000000000000001010100110011", -- 5426 FREE #<CONS 0 5427>
 "00000000000000000001010100110100", -- 5427 FREE #<CONS 0 5428>
 "00000000000000000001010100110101", -- 5428 FREE #<CONS 0 5429>
 "00000000000000000001010100110110", -- 5429 FREE #<CONS 0 5430>
 "00000000000000000001010100110111", -- 5430 FREE #<CONS 0 5431>
 "00000000000000000001010100111000", -- 5431 FREE #<CONS 0 5432>
 "00000000000000000001010100111001", -- 5432 FREE #<CONS 0 5433>
 "00000000000000000001010100111010", -- 5433 FREE #<CONS 0 5434>
 "00000000000000000001010100111011", -- 5434 FREE #<CONS 0 5435>
 "00000000000000000001010100111100", -- 5435 FREE #<CONS 0 5436>
 "00000000000000000001010100111101", -- 5436 FREE #<CONS 0 5437>
 "00000000000000000001010100111110", -- 5437 FREE #<CONS 0 5438>
 "00000000000000000001010100111111", -- 5438 FREE #<CONS 0 5439>
 "00000000000000000001010101000000", -- 5439 FREE #<CONS 0 5440>
 "00000000000000000001010101000001", -- 5440 FREE #<CONS 0 5441>
 "00000000000000000001010101000010", -- 5441 FREE #<CONS 0 5442>
 "00000000000000000001010101000011", -- 5442 FREE #<CONS 0 5443>
 "00000000000000000001010101000100", -- 5443 FREE #<CONS 0 5444>
 "00000000000000000001010101000101", -- 5444 FREE #<CONS 0 5445>
 "00000000000000000001010101000110", -- 5445 FREE #<CONS 0 5446>
 "00000000000000000001010101000111", -- 5446 FREE #<CONS 0 5447>
 "00000000000000000001010101001000", -- 5447 FREE #<CONS 0 5448>
 "00000000000000000001010101001001", -- 5448 FREE #<CONS 0 5449>
 "00000000000000000001010101001010", -- 5449 FREE #<CONS 0 5450>
 "00000000000000000001010101001011", -- 5450 FREE #<CONS 0 5451>
 "00000000000000000001010101001100", -- 5451 FREE #<CONS 0 5452>
 "00000000000000000001010101001101", -- 5452 FREE #<CONS 0 5453>
 "00000000000000000001010101001110", -- 5453 FREE #<CONS 0 5454>
 "00000000000000000001010101001111", -- 5454 FREE #<CONS 0 5455>
 "00000000000000000001010101010000", -- 5455 FREE #<CONS 0 5456>
 "00000000000000000001010101010001", -- 5456 FREE #<CONS 0 5457>
 "00000000000000000001010101010010", -- 5457 FREE #<CONS 0 5458>
 "00000000000000000001010101010011", -- 5458 FREE #<CONS 0 5459>
 "00000000000000000001010101010100", -- 5459 FREE #<CONS 0 5460>
 "00000000000000000001010101010101", -- 5460 FREE #<CONS 0 5461>
 "00000000000000000001010101010110", -- 5461 FREE #<CONS 0 5462>
 "00000000000000000001010101010111", -- 5462 FREE #<CONS 0 5463>
 "00000000000000000001010101011000", -- 5463 FREE #<CONS 0 5464>
 "00000000000000000001010101011001", -- 5464 FREE #<CONS 0 5465>
 "00000000000000000001010101011010", -- 5465 FREE #<CONS 0 5466>
 "00000000000000000001010101011011", -- 5466 FREE #<CONS 0 5467>
 "00000000000000000001010101011100", -- 5467 FREE #<CONS 0 5468>
 "00000000000000000001010101011101", -- 5468 FREE #<CONS 0 5469>
 "00000000000000000001010101011110", -- 5469 FREE #<CONS 0 5470>
 "00000000000000000001010101011111", -- 5470 FREE #<CONS 0 5471>
 "00000000000000000001010101100000", -- 5471 FREE #<CONS 0 5472>
 "00000000000000000001010101100001", -- 5472 FREE #<CONS 0 5473>
 "00000000000000000001010101100010", -- 5473 FREE #<CONS 0 5474>
 "00000000000000000001010101100011", -- 5474 FREE #<CONS 0 5475>
 "00000000000000000001010101100100", -- 5475 FREE #<CONS 0 5476>
 "00000000000000000001010101100101", -- 5476 FREE #<CONS 0 5477>
 "00000000000000000001010101100110", -- 5477 FREE #<CONS 0 5478>
 "00000000000000000001010101100111", -- 5478 FREE #<CONS 0 5479>
 "00000000000000000001010101101000", -- 5479 FREE #<CONS 0 5480>
 "00000000000000000001010101101001", -- 5480 FREE #<CONS 0 5481>
 "00000000000000000001010101101010", -- 5481 FREE #<CONS 0 5482>
 "00000000000000000001010101101011", -- 5482 FREE #<CONS 0 5483>
 "00000000000000000001010101101100", -- 5483 FREE #<CONS 0 5484>
 "00000000000000000001010101101101", -- 5484 FREE #<CONS 0 5485>
 "00000000000000000001010101101110", -- 5485 FREE #<CONS 0 5486>
 "00000000000000000001010101101111", -- 5486 FREE #<CONS 0 5487>
 "00000000000000000001010101110000", -- 5487 FREE #<CONS 0 5488>
 "00000000000000000001010101110001", -- 5488 FREE #<CONS 0 5489>
 "00000000000000000001010101110010", -- 5489 FREE #<CONS 0 5490>
 "00000000000000000001010101110011", -- 5490 FREE #<CONS 0 5491>
 "00000000000000000001010101110100", -- 5491 FREE #<CONS 0 5492>
 "00000000000000000001010101110101", -- 5492 FREE #<CONS 0 5493>
 "00000000000000000001010101110110", -- 5493 FREE #<CONS 0 5494>
 "00000000000000000001010101110111", -- 5494 FREE #<CONS 0 5495>
 "00000000000000000001010101111000", -- 5495 FREE #<CONS 0 5496>
 "00000000000000000001010101111001", -- 5496 FREE #<CONS 0 5497>
 "00000000000000000001010101111010", -- 5497 FREE #<CONS 0 5498>
 "00000000000000000001010101111011", -- 5498 FREE #<CONS 0 5499>
 "00000000000000000001010101111100", -- 5499 FREE #<CONS 0 5500>
 "00000000000000000001010101111101", -- 5500 FREE #<CONS 0 5501>
 "00000000000000000001010101111110", -- 5501 FREE #<CONS 0 5502>
 "00000000000000000001010101111111", -- 5502 FREE #<CONS 0 5503>
 "00000000000000000001010110000000", -- 5503 FREE #<CONS 0 5504>
 "00000000000000000001010110000001", -- 5504 FREE #<CONS 0 5505>
 "00000000000000000001010110000010", -- 5505 FREE #<CONS 0 5506>
 "00000000000000000001010110000011", -- 5506 FREE #<CONS 0 5507>
 "00000000000000000001010110000100", -- 5507 FREE #<CONS 0 5508>
 "00000000000000000001010110000101", -- 5508 FREE #<CONS 0 5509>
 "00000000000000000001010110000110", -- 5509 FREE #<CONS 0 5510>
 "00000000000000000001010110000111", -- 5510 FREE #<CONS 0 5511>
 "00000000000000000001010110001000", -- 5511 FREE #<CONS 0 5512>
 "00000000000000000001010110001001", -- 5512 FREE #<CONS 0 5513>
 "00000000000000000001010110001010", -- 5513 FREE #<CONS 0 5514>
 "00000000000000000001010110001011", -- 5514 FREE #<CONS 0 5515>
 "00000000000000000001010110001100", -- 5515 FREE #<CONS 0 5516>
 "00000000000000000001010110001101", -- 5516 FREE #<CONS 0 5517>
 "00000000000000000001010110001110", -- 5517 FREE #<CONS 0 5518>
 "00000000000000000001010110001111", -- 5518 FREE #<CONS 0 5519>
 "00000000000000000001010110010000", -- 5519 FREE #<CONS 0 5520>
 "00000000000000000001010110010001", -- 5520 FREE #<CONS 0 5521>
 "00000000000000000001010110010010", -- 5521 FREE #<CONS 0 5522>
 "00000000000000000001010110010011", -- 5522 FREE #<CONS 0 5523>
 "00000000000000000001010110010100", -- 5523 FREE #<CONS 0 5524>
 "00000000000000000001010110010101", -- 5524 FREE #<CONS 0 5525>
 "00000000000000000001010110010110", -- 5525 FREE #<CONS 0 5526>
 "00000000000000000001010110010111", -- 5526 FREE #<CONS 0 5527>
 "00000000000000000001010110011000", -- 5527 FREE #<CONS 0 5528>
 "00000000000000000001010110011001", -- 5528 FREE #<CONS 0 5529>
 "00000000000000000001010110011010", -- 5529 FREE #<CONS 0 5530>
 "00000000000000000001010110011011", -- 5530 FREE #<CONS 0 5531>
 "00000000000000000001010110011100", -- 5531 FREE #<CONS 0 5532>
 "00000000000000000001010110011101", -- 5532 FREE #<CONS 0 5533>
 "00000000000000000001010110011110", -- 5533 FREE #<CONS 0 5534>
 "00000000000000000001010110011111", -- 5534 FREE #<CONS 0 5535>
 "00000000000000000001010110100000", -- 5535 FREE #<CONS 0 5536>
 "00000000000000000001010110100001", -- 5536 FREE #<CONS 0 5537>
 "00000000000000000001010110100010", -- 5537 FREE #<CONS 0 5538>
 "00000000000000000001010110100011", -- 5538 FREE #<CONS 0 5539>
 "00000000000000000001010110100100", -- 5539 FREE #<CONS 0 5540>
 "00000000000000000001010110100101", -- 5540 FREE #<CONS 0 5541>
 "00000000000000000001010110100110", -- 5541 FREE #<CONS 0 5542>
 "00000000000000000001010110100111", -- 5542 FREE #<CONS 0 5543>
 "00000000000000000001010110101000", -- 5543 FREE #<CONS 0 5544>
 "00000000000000000001010110101001", -- 5544 FREE #<CONS 0 5545>
 "00000000000000000001010110101010", -- 5545 FREE #<CONS 0 5546>
 "00000000000000000001010110101011", -- 5546 FREE #<CONS 0 5547>
 "00000000000000000001010110101100", -- 5547 FREE #<CONS 0 5548>
 "00000000000000000001010110101101", -- 5548 FREE #<CONS 0 5549>
 "00000000000000000001010110101110", -- 5549 FREE #<CONS 0 5550>
 "00000000000000000001010110101111", -- 5550 FREE #<CONS 0 5551>
 "00000000000000000001010110110000", -- 5551 FREE #<CONS 0 5552>
 "00000000000000000001010110110001", -- 5552 FREE #<CONS 0 5553>
 "00000000000000000001010110110010", -- 5553 FREE #<CONS 0 5554>
 "00000000000000000001010110110011", -- 5554 FREE #<CONS 0 5555>
 "00000000000000000001010110110100", -- 5555 FREE #<CONS 0 5556>
 "00000000000000000001010110110101", -- 5556 FREE #<CONS 0 5557>
 "00000000000000000001010110110110", -- 5557 FREE #<CONS 0 5558>
 "00000000000000000001010110110111", -- 5558 FREE #<CONS 0 5559>
 "00000000000000000001010110111000", -- 5559 FREE #<CONS 0 5560>
 "00000000000000000001010110111001", -- 5560 FREE #<CONS 0 5561>
 "00000000000000000001010110111010", -- 5561 FREE #<CONS 0 5562>
 "00000000000000000001010110111011", -- 5562 FREE #<CONS 0 5563>
 "00000000000000000001010110111100", -- 5563 FREE #<CONS 0 5564>
 "00000000000000000001010110111101", -- 5564 FREE #<CONS 0 5565>
 "00000000000000000001010110111110", -- 5565 FREE #<CONS 0 5566>
 "00000000000000000001010110111111", -- 5566 FREE #<CONS 0 5567>
 "00000000000000000001010111000000", -- 5567 FREE #<CONS 0 5568>
 "00000000000000000001010111000001", -- 5568 FREE #<CONS 0 5569>
 "00000000000000000001010111000010", -- 5569 FREE #<CONS 0 5570>
 "00000000000000000001010111000011", -- 5570 FREE #<CONS 0 5571>
 "00000000000000000001010111000100", -- 5571 FREE #<CONS 0 5572>
 "00000000000000000001010111000101", -- 5572 FREE #<CONS 0 5573>
 "00000000000000000001010111000110", -- 5573 FREE #<CONS 0 5574>
 "00000000000000000001010111000111", -- 5574 FREE #<CONS 0 5575>
 "00000000000000000001010111001000", -- 5575 FREE #<CONS 0 5576>
 "00000000000000000001010111001001", -- 5576 FREE #<CONS 0 5577>
 "00000000000000000001010111001010", -- 5577 FREE #<CONS 0 5578>
 "00000000000000000001010111001011", -- 5578 FREE #<CONS 0 5579>
 "00000000000000000001010111001100", -- 5579 FREE #<CONS 0 5580>
 "00000000000000000001010111001101", -- 5580 FREE #<CONS 0 5581>
 "00000000000000000001010111001110", -- 5581 FREE #<CONS 0 5582>
 "00000000000000000001010111001111", -- 5582 FREE #<CONS 0 5583>
 "00000000000000000001010111010000", -- 5583 FREE #<CONS 0 5584>
 "00000000000000000001010111010001", -- 5584 FREE #<CONS 0 5585>
 "00000000000000000001010111010010", -- 5585 FREE #<CONS 0 5586>
 "00000000000000000001010111010011", -- 5586 FREE #<CONS 0 5587>
 "00000000000000000001010111010100", -- 5587 FREE #<CONS 0 5588>
 "00000000000000000001010111010101", -- 5588 FREE #<CONS 0 5589>
 "00000000000000000001010111010110", -- 5589 FREE #<CONS 0 5590>
 "00000000000000000001010111010111", -- 5590 FREE #<CONS 0 5591>
 "00000000000000000001010111011000", -- 5591 FREE #<CONS 0 5592>
 "00000000000000000001010111011001", -- 5592 FREE #<CONS 0 5593>
 "00000000000000000001010111011010", -- 5593 FREE #<CONS 0 5594>
 "00000000000000000001010111011011", -- 5594 FREE #<CONS 0 5595>
 "00000000000000000001010111011100", -- 5595 FREE #<CONS 0 5596>
 "00000000000000000001010111011101", -- 5596 FREE #<CONS 0 5597>
 "00000000000000000001010111011110", -- 5597 FREE #<CONS 0 5598>
 "00000000000000000001010111011111", -- 5598 FREE #<CONS 0 5599>
 "00000000000000000001010111100000", -- 5599 FREE #<CONS 0 5600>
 "00000000000000000001010111100001", -- 5600 FREE #<CONS 0 5601>
 "00000000000000000001010111100010", -- 5601 FREE #<CONS 0 5602>
 "00000000000000000001010111100011", -- 5602 FREE #<CONS 0 5603>
 "00000000000000000001010111100100", -- 5603 FREE #<CONS 0 5604>
 "00000000000000000001010111100101", -- 5604 FREE #<CONS 0 5605>
 "00000000000000000001010111100110", -- 5605 FREE #<CONS 0 5606>
 "00000000000000000001010111100111", -- 5606 FREE #<CONS 0 5607>
 "00000000000000000001010111101000", -- 5607 FREE #<CONS 0 5608>
 "00000000000000000001010111101001", -- 5608 FREE #<CONS 0 5609>
 "00000000000000000001010111101010", -- 5609 FREE #<CONS 0 5610>
 "00000000000000000001010111101011", -- 5610 FREE #<CONS 0 5611>
 "00000000000000000001010111101100", -- 5611 FREE #<CONS 0 5612>
 "00000000000000000001010111101101", -- 5612 FREE #<CONS 0 5613>
 "00000000000000000001010111101110", -- 5613 FREE #<CONS 0 5614>
 "00000000000000000001010111101111", -- 5614 FREE #<CONS 0 5615>
 "00000000000000000001010111110000", -- 5615 FREE #<CONS 0 5616>
 "00000000000000000001010111110001", -- 5616 FREE #<CONS 0 5617>
 "00000000000000000001010111110010", -- 5617 FREE #<CONS 0 5618>
 "00000000000000000001010111110011", -- 5618 FREE #<CONS 0 5619>
 "00000000000000000001010111110100", -- 5619 FREE #<CONS 0 5620>
 "00000000000000000001010111110101", -- 5620 FREE #<CONS 0 5621>
 "00000000000000000001010111110110", -- 5621 FREE #<CONS 0 5622>
 "00000000000000000001010111110111", -- 5622 FREE #<CONS 0 5623>
 "00000000000000000001010111111000", -- 5623 FREE #<CONS 0 5624>
 "00000000000000000001010111111001", -- 5624 FREE #<CONS 0 5625>
 "00000000000000000001010111111010", -- 5625 FREE #<CONS 0 5626>
 "00000000000000000001010111111011", -- 5626 FREE #<CONS 0 5627>
 "00000000000000000001010111111100", -- 5627 FREE #<CONS 0 5628>
 "00000000000000000001010111111101", -- 5628 FREE #<CONS 0 5629>
 "00000000000000000001010111111110", -- 5629 FREE #<CONS 0 5630>
 "00000000000000000001010111111111", -- 5630 FREE #<CONS 0 5631>
 "00000000000000000001011000000000", -- 5631 FREE #<CONS 0 5632>
 "00000000000000000001011000000001", -- 5632 FREE #<CONS 0 5633>
 "00000000000000000001011000000010", -- 5633 FREE #<CONS 0 5634>
 "00000000000000000001011000000011", -- 5634 FREE #<CONS 0 5635>
 "00000000000000000001011000000100", -- 5635 FREE #<CONS 0 5636>
 "00000000000000000001011000000101", -- 5636 FREE #<CONS 0 5637>
 "00000000000000000001011000000110", -- 5637 FREE #<CONS 0 5638>
 "00000000000000000001011000000111", -- 5638 FREE #<CONS 0 5639>
 "00000000000000000001011000001000", -- 5639 FREE #<CONS 0 5640>
 "00000000000000000001011000001001", -- 5640 FREE #<CONS 0 5641>
 "00000000000000000001011000001010", -- 5641 FREE #<CONS 0 5642>
 "00000000000000000001011000001011", -- 5642 FREE #<CONS 0 5643>
 "00000000000000000001011000001100", -- 5643 FREE #<CONS 0 5644>
 "00000000000000000001011000001101", -- 5644 FREE #<CONS 0 5645>
 "00000000000000000001011000001110", -- 5645 FREE #<CONS 0 5646>
 "00000000000000000001011000001111", -- 5646 FREE #<CONS 0 5647>
 "00000000000000000001011000010000", -- 5647 FREE #<CONS 0 5648>
 "00000000000000000001011000010001", -- 5648 FREE #<CONS 0 5649>
 "00000000000000000001011000010010", -- 5649 FREE #<CONS 0 5650>
 "00000000000000000001011000010011", -- 5650 FREE #<CONS 0 5651>
 "00000000000000000001011000010100", -- 5651 FREE #<CONS 0 5652>
 "00000000000000000001011000010101", -- 5652 FREE #<CONS 0 5653>
 "00000000000000000001011000010110", -- 5653 FREE #<CONS 0 5654>
 "00000000000000000001011000010111", -- 5654 FREE #<CONS 0 5655>
 "00000000000000000001011000011000", -- 5655 FREE #<CONS 0 5656>
 "00000000000000000001011000011001", -- 5656 FREE #<CONS 0 5657>
 "00000000000000000001011000011010", -- 5657 FREE #<CONS 0 5658>
 "00000000000000000001011000011011", -- 5658 FREE #<CONS 0 5659>
 "00000000000000000001011000011100", -- 5659 FREE #<CONS 0 5660>
 "00000000000000000001011000011101", -- 5660 FREE #<CONS 0 5661>
 "00000000000000000001011000011110", -- 5661 FREE #<CONS 0 5662>
 "00000000000000000001011000011111", -- 5662 FREE #<CONS 0 5663>
 "00000000000000000001011000100000", -- 5663 FREE #<CONS 0 5664>
 "00000000000000000001011000100001", -- 5664 FREE #<CONS 0 5665>
 "00000000000000000001011000100010", -- 5665 FREE #<CONS 0 5666>
 "00000000000000000001011000100011", -- 5666 FREE #<CONS 0 5667>
 "00000000000000000001011000100100", -- 5667 FREE #<CONS 0 5668>
 "00000000000000000001011000100101", -- 5668 FREE #<CONS 0 5669>
 "00000000000000000001011000100110", -- 5669 FREE #<CONS 0 5670>
 "00000000000000000001011000100111", -- 5670 FREE #<CONS 0 5671>
 "00000000000000000001011000101000", -- 5671 FREE #<CONS 0 5672>
 "00000000000000000001011000101001", -- 5672 FREE #<CONS 0 5673>
 "00000000000000000001011000101010", -- 5673 FREE #<CONS 0 5674>
 "00000000000000000001011000101011", -- 5674 FREE #<CONS 0 5675>
 "00000000000000000001011000101100", -- 5675 FREE #<CONS 0 5676>
 "00000000000000000001011000101101", -- 5676 FREE #<CONS 0 5677>
 "00000000000000000001011000101110", -- 5677 FREE #<CONS 0 5678>
 "00000000000000000001011000101111", -- 5678 FREE #<CONS 0 5679>
 "00000000000000000001011000110000", -- 5679 FREE #<CONS 0 5680>
 "00000000000000000001011000110001", -- 5680 FREE #<CONS 0 5681>
 "00000000000000000001011000110010", -- 5681 FREE #<CONS 0 5682>
 "00000000000000000001011000110011", -- 5682 FREE #<CONS 0 5683>
 "00000000000000000001011000110100", -- 5683 FREE #<CONS 0 5684>
 "00000000000000000001011000110101", -- 5684 FREE #<CONS 0 5685>
 "00000000000000000001011000110110", -- 5685 FREE #<CONS 0 5686>
 "00000000000000000001011000110111", -- 5686 FREE #<CONS 0 5687>
 "00000000000000000001011000111000", -- 5687 FREE #<CONS 0 5688>
 "00000000000000000001011000111001", -- 5688 FREE #<CONS 0 5689>
 "00000000000000000001011000111010", -- 5689 FREE #<CONS 0 5690>
 "00000000000000000001011000111011", -- 5690 FREE #<CONS 0 5691>
 "00000000000000000001011000111100", -- 5691 FREE #<CONS 0 5692>
 "00000000000000000001011000111101", -- 5692 FREE #<CONS 0 5693>
 "00000000000000000001011000111110", -- 5693 FREE #<CONS 0 5694>
 "00000000000000000001011000111111", -- 5694 FREE #<CONS 0 5695>
 "00000000000000000001011001000000", -- 5695 FREE #<CONS 0 5696>
 "00000000000000000001011001000001", -- 5696 FREE #<CONS 0 5697>
 "00000000000000000001011001000010", -- 5697 FREE #<CONS 0 5698>
 "00000000000000000001011001000011", -- 5698 FREE #<CONS 0 5699>
 "00000000000000000001011001000100", -- 5699 FREE #<CONS 0 5700>
 "00000000000000000001011001000101", -- 5700 FREE #<CONS 0 5701>
 "00000000000000000001011001000110", -- 5701 FREE #<CONS 0 5702>
 "00000000000000000001011001000111", -- 5702 FREE #<CONS 0 5703>
 "00000000000000000001011001001000", -- 5703 FREE #<CONS 0 5704>
 "00000000000000000001011001001001", -- 5704 FREE #<CONS 0 5705>
 "00000000000000000001011001001010", -- 5705 FREE #<CONS 0 5706>
 "00000000000000000001011001001011", -- 5706 FREE #<CONS 0 5707>
 "00000000000000000001011001001100", -- 5707 FREE #<CONS 0 5708>
 "00000000000000000001011001001101", -- 5708 FREE #<CONS 0 5709>
 "00000000000000000001011001001110", -- 5709 FREE #<CONS 0 5710>
 "00000000000000000001011001001111", -- 5710 FREE #<CONS 0 5711>
 "00000000000000000001011001010000", -- 5711 FREE #<CONS 0 5712>
 "00000000000000000001011001010001", -- 5712 FREE #<CONS 0 5713>
 "00000000000000000001011001010010", -- 5713 FREE #<CONS 0 5714>
 "00000000000000000001011001010011", -- 5714 FREE #<CONS 0 5715>
 "00000000000000000001011001010100", -- 5715 FREE #<CONS 0 5716>
 "00000000000000000001011001010101", -- 5716 FREE #<CONS 0 5717>
 "00000000000000000001011001010110", -- 5717 FREE #<CONS 0 5718>
 "00000000000000000001011001010111", -- 5718 FREE #<CONS 0 5719>
 "00000000000000000001011001011000", -- 5719 FREE #<CONS 0 5720>
 "00000000000000000001011001011001", -- 5720 FREE #<CONS 0 5721>
 "00000000000000000001011001011010", -- 5721 FREE #<CONS 0 5722>
 "00000000000000000001011001011011", -- 5722 FREE #<CONS 0 5723>
 "00000000000000000001011001011100", -- 5723 FREE #<CONS 0 5724>
 "00000000000000000001011001011101", -- 5724 FREE #<CONS 0 5725>
 "00000000000000000001011001011110", -- 5725 FREE #<CONS 0 5726>
 "00000000000000000001011001011111", -- 5726 FREE #<CONS 0 5727>
 "00000000000000000001011001100000", -- 5727 FREE #<CONS 0 5728>
 "00000000000000000001011001100001", -- 5728 FREE #<CONS 0 5729>
 "00000000000000000001011001100010", -- 5729 FREE #<CONS 0 5730>
 "00000000000000000001011001100011", -- 5730 FREE #<CONS 0 5731>
 "00000000000000000001011001100100", -- 5731 FREE #<CONS 0 5732>
 "00000000000000000001011001100101", -- 5732 FREE #<CONS 0 5733>
 "00000000000000000001011001100110", -- 5733 FREE #<CONS 0 5734>
 "00000000000000000001011001100111", -- 5734 FREE #<CONS 0 5735>
 "00000000000000000001011001101000", -- 5735 FREE #<CONS 0 5736>
 "00000000000000000001011001101001", -- 5736 FREE #<CONS 0 5737>
 "00000000000000000001011001101010", -- 5737 FREE #<CONS 0 5738>
 "00000000000000000001011001101011", -- 5738 FREE #<CONS 0 5739>
 "00000000000000000001011001101100", -- 5739 FREE #<CONS 0 5740>
 "00000000000000000001011001101101", -- 5740 FREE #<CONS 0 5741>
 "00000000000000000001011001101110", -- 5741 FREE #<CONS 0 5742>
 "00000000000000000001011001101111", -- 5742 FREE #<CONS 0 5743>
 "00000000000000000001011001110000", -- 5743 FREE #<CONS 0 5744>
 "00000000000000000001011001110001", -- 5744 FREE #<CONS 0 5745>
 "00000000000000000001011001110010", -- 5745 FREE #<CONS 0 5746>
 "00000000000000000001011001110011", -- 5746 FREE #<CONS 0 5747>
 "00000000000000000001011001110100", -- 5747 FREE #<CONS 0 5748>
 "00000000000000000001011001110101", -- 5748 FREE #<CONS 0 5749>
 "00000000000000000001011001110110", -- 5749 FREE #<CONS 0 5750>
 "00000000000000000001011001110111", -- 5750 FREE #<CONS 0 5751>
 "00000000000000000001011001111000", -- 5751 FREE #<CONS 0 5752>
 "00000000000000000001011001111001", -- 5752 FREE #<CONS 0 5753>
 "00000000000000000001011001111010", -- 5753 FREE #<CONS 0 5754>
 "00000000000000000001011001111011", -- 5754 FREE #<CONS 0 5755>
 "00000000000000000001011001111100", -- 5755 FREE #<CONS 0 5756>
 "00000000000000000001011001111101", -- 5756 FREE #<CONS 0 5757>
 "00000000000000000001011001111110", -- 5757 FREE #<CONS 0 5758>
 "00000000000000000001011001111111", -- 5758 FREE #<CONS 0 5759>
 "00000000000000000001011010000000", -- 5759 FREE #<CONS 0 5760>
 "00000000000000000001011010000001", -- 5760 FREE #<CONS 0 5761>
 "00000000000000000001011010000010", -- 5761 FREE #<CONS 0 5762>
 "00000000000000000001011010000011", -- 5762 FREE #<CONS 0 5763>
 "00000000000000000001011010000100", -- 5763 FREE #<CONS 0 5764>
 "00000000000000000001011010000101", -- 5764 FREE #<CONS 0 5765>
 "00000000000000000001011010000110", -- 5765 FREE #<CONS 0 5766>
 "00000000000000000001011010000111", -- 5766 FREE #<CONS 0 5767>
 "00000000000000000001011010001000", -- 5767 FREE #<CONS 0 5768>
 "00000000000000000001011010001001", -- 5768 FREE #<CONS 0 5769>
 "00000000000000000001011010001010", -- 5769 FREE #<CONS 0 5770>
 "00000000000000000001011010001011", -- 5770 FREE #<CONS 0 5771>
 "00000000000000000001011010001100", -- 5771 FREE #<CONS 0 5772>
 "00000000000000000001011010001101", -- 5772 FREE #<CONS 0 5773>
 "00000000000000000001011010001110", -- 5773 FREE #<CONS 0 5774>
 "00000000000000000001011010001111", -- 5774 FREE #<CONS 0 5775>
 "00000000000000000001011010010000", -- 5775 FREE #<CONS 0 5776>
 "00000000000000000001011010010001", -- 5776 FREE #<CONS 0 5777>
 "00000000000000000001011010010010", -- 5777 FREE #<CONS 0 5778>
 "00000000000000000001011010010011", -- 5778 FREE #<CONS 0 5779>
 "00000000000000000001011010010100", -- 5779 FREE #<CONS 0 5780>
 "00000000000000000001011010010101", -- 5780 FREE #<CONS 0 5781>
 "00000000000000000001011010010110", -- 5781 FREE #<CONS 0 5782>
 "00000000000000000001011010010111", -- 5782 FREE #<CONS 0 5783>
 "00000000000000000001011010011000", -- 5783 FREE #<CONS 0 5784>
 "00000000000000000001011010011001", -- 5784 FREE #<CONS 0 5785>
 "00000000000000000001011010011010", -- 5785 FREE #<CONS 0 5786>
 "00000000000000000001011010011011", -- 5786 FREE #<CONS 0 5787>
 "00000000000000000001011010011100", -- 5787 FREE #<CONS 0 5788>
 "00000000000000000001011010011101", -- 5788 FREE #<CONS 0 5789>
 "00000000000000000001011010011110", -- 5789 FREE #<CONS 0 5790>
 "00000000000000000001011010011111", -- 5790 FREE #<CONS 0 5791>
 "00000000000000000001011010100000", -- 5791 FREE #<CONS 0 5792>
 "00000000000000000001011010100001", -- 5792 FREE #<CONS 0 5793>
 "00000000000000000001011010100010", -- 5793 FREE #<CONS 0 5794>
 "00000000000000000001011010100011", -- 5794 FREE #<CONS 0 5795>
 "00000000000000000001011010100100", -- 5795 FREE #<CONS 0 5796>
 "00000000000000000001011010100101", -- 5796 FREE #<CONS 0 5797>
 "00000000000000000001011010100110", -- 5797 FREE #<CONS 0 5798>
 "00000000000000000001011010100111", -- 5798 FREE #<CONS 0 5799>
 "00000000000000000001011010101000", -- 5799 FREE #<CONS 0 5800>
 "00000000000000000001011010101001", -- 5800 FREE #<CONS 0 5801>
 "00000000000000000001011010101010", -- 5801 FREE #<CONS 0 5802>
 "00000000000000000001011010101011", -- 5802 FREE #<CONS 0 5803>
 "00000000000000000001011010101100", -- 5803 FREE #<CONS 0 5804>
 "00000000000000000001011010101101", -- 5804 FREE #<CONS 0 5805>
 "00000000000000000001011010101110", -- 5805 FREE #<CONS 0 5806>
 "00000000000000000001011010101111", -- 5806 FREE #<CONS 0 5807>
 "00000000000000000001011010110000", -- 5807 FREE #<CONS 0 5808>
 "00000000000000000001011010110001", -- 5808 FREE #<CONS 0 5809>
 "00000000000000000001011010110010", -- 5809 FREE #<CONS 0 5810>
 "00000000000000000001011010110011", -- 5810 FREE #<CONS 0 5811>
 "00000000000000000001011010110100", -- 5811 FREE #<CONS 0 5812>
 "00000000000000000001011010110101", -- 5812 FREE #<CONS 0 5813>
 "00000000000000000001011010110110", -- 5813 FREE #<CONS 0 5814>
 "00000000000000000001011010110111", -- 5814 FREE #<CONS 0 5815>
 "00000000000000000001011010111000", -- 5815 FREE #<CONS 0 5816>
 "00000000000000000001011010111001", -- 5816 FREE #<CONS 0 5817>
 "00000000000000000001011010111010", -- 5817 FREE #<CONS 0 5818>
 "00000000000000000001011010111011", -- 5818 FREE #<CONS 0 5819>
 "00000000000000000001011010111100", -- 5819 FREE #<CONS 0 5820>
 "00000000000000000001011010111101", -- 5820 FREE #<CONS 0 5821>
 "00000000000000000001011010111110", -- 5821 FREE #<CONS 0 5822>
 "00000000000000000001011010111111", -- 5822 FREE #<CONS 0 5823>
 "00000000000000000001011011000000", -- 5823 FREE #<CONS 0 5824>
 "00000000000000000001011011000001", -- 5824 FREE #<CONS 0 5825>
 "00000000000000000001011011000010", -- 5825 FREE #<CONS 0 5826>
 "00000000000000000001011011000011", -- 5826 FREE #<CONS 0 5827>
 "00000000000000000001011011000100", -- 5827 FREE #<CONS 0 5828>
 "00000000000000000001011011000101", -- 5828 FREE #<CONS 0 5829>
 "00000000000000000001011011000110", -- 5829 FREE #<CONS 0 5830>
 "00000000000000000001011011000111", -- 5830 FREE #<CONS 0 5831>
 "00000000000000000001011011001000", -- 5831 FREE #<CONS 0 5832>
 "00000000000000000001011011001001", -- 5832 FREE #<CONS 0 5833>
 "00000000000000000001011011001010", -- 5833 FREE #<CONS 0 5834>
 "00000000000000000001011011001011", -- 5834 FREE #<CONS 0 5835>
 "00000000000000000001011011001100", -- 5835 FREE #<CONS 0 5836>
 "00000000000000000001011011001101", -- 5836 FREE #<CONS 0 5837>
 "00000000000000000001011011001110", -- 5837 FREE #<CONS 0 5838>
 "00000000000000000001011011001111", -- 5838 FREE #<CONS 0 5839>
 "00000000000000000001011011010000", -- 5839 FREE #<CONS 0 5840>
 "00000000000000000001011011010001", -- 5840 FREE #<CONS 0 5841>
 "00000000000000000001011011010010", -- 5841 FREE #<CONS 0 5842>
 "00000000000000000001011011010011", -- 5842 FREE #<CONS 0 5843>
 "00000000000000000001011011010100", -- 5843 FREE #<CONS 0 5844>
 "00000000000000000001011011010101", -- 5844 FREE #<CONS 0 5845>
 "00000000000000000001011011010110", -- 5845 FREE #<CONS 0 5846>
 "00000000000000000001011011010111", -- 5846 FREE #<CONS 0 5847>
 "00000000000000000001011011011000", -- 5847 FREE #<CONS 0 5848>
 "00000000000000000001011011011001", -- 5848 FREE #<CONS 0 5849>
 "00000000000000000001011011011010", -- 5849 FREE #<CONS 0 5850>
 "00000000000000000001011011011011", -- 5850 FREE #<CONS 0 5851>
 "00000000000000000001011011011100", -- 5851 FREE #<CONS 0 5852>
 "00000000000000000001011011011101", -- 5852 FREE #<CONS 0 5853>
 "00000000000000000001011011011110", -- 5853 FREE #<CONS 0 5854>
 "00000000000000000001011011011111", -- 5854 FREE #<CONS 0 5855>
 "00000000000000000001011011100000", -- 5855 FREE #<CONS 0 5856>
 "00000000000000000001011011100001", -- 5856 FREE #<CONS 0 5857>
 "00000000000000000001011011100010", -- 5857 FREE #<CONS 0 5858>
 "00000000000000000001011011100011", -- 5858 FREE #<CONS 0 5859>
 "00000000000000000001011011100100", -- 5859 FREE #<CONS 0 5860>
 "00000000000000000001011011100101", -- 5860 FREE #<CONS 0 5861>
 "00000000000000000001011011100110", -- 5861 FREE #<CONS 0 5862>
 "00000000000000000001011011100111", -- 5862 FREE #<CONS 0 5863>
 "00000000000000000001011011101000", -- 5863 FREE #<CONS 0 5864>
 "00000000000000000001011011101001", -- 5864 FREE #<CONS 0 5865>
 "00000000000000000001011011101010", -- 5865 FREE #<CONS 0 5866>
 "00000000000000000001011011101011", -- 5866 FREE #<CONS 0 5867>
 "00000000000000000001011011101100", -- 5867 FREE #<CONS 0 5868>
 "00000000000000000001011011101101", -- 5868 FREE #<CONS 0 5869>
 "00000000000000000001011011101110", -- 5869 FREE #<CONS 0 5870>
 "00000000000000000001011011101111", -- 5870 FREE #<CONS 0 5871>
 "00000000000000000001011011110000", -- 5871 FREE #<CONS 0 5872>
 "00000000000000000001011011110001", -- 5872 FREE #<CONS 0 5873>
 "00000000000000000001011011110010", -- 5873 FREE #<CONS 0 5874>
 "00000000000000000001011011110011", -- 5874 FREE #<CONS 0 5875>
 "00000000000000000001011011110100", -- 5875 FREE #<CONS 0 5876>
 "00000000000000000001011011110101", -- 5876 FREE #<CONS 0 5877>
 "00000000000000000001011011110110", -- 5877 FREE #<CONS 0 5878>
 "00000000000000000001011011110111", -- 5878 FREE #<CONS 0 5879>
 "00000000000000000001011011111000", -- 5879 FREE #<CONS 0 5880>
 "00000000000000000001011011111001", -- 5880 FREE #<CONS 0 5881>
 "00000000000000000001011011111010", -- 5881 FREE #<CONS 0 5882>
 "00000000000000000001011011111011", -- 5882 FREE #<CONS 0 5883>
 "00000000000000000001011011111100", -- 5883 FREE #<CONS 0 5884>
 "00000000000000000001011011111101", -- 5884 FREE #<CONS 0 5885>
 "00000000000000000001011011111110", -- 5885 FREE #<CONS 0 5886>
 "00000000000000000001011011111111", -- 5886 FREE #<CONS 0 5887>
 "00000000000000000001011100000000", -- 5887 FREE #<CONS 0 5888>
 "00000000000000000001011100000001", -- 5888 FREE #<CONS 0 5889>
 "00000000000000000001011100000010", -- 5889 FREE #<CONS 0 5890>
 "00000000000000000001011100000011", -- 5890 FREE #<CONS 0 5891>
 "00000000000000000001011100000100", -- 5891 FREE #<CONS 0 5892>
 "00000000000000000001011100000101", -- 5892 FREE #<CONS 0 5893>
 "00000000000000000001011100000110", -- 5893 FREE #<CONS 0 5894>
 "00000000000000000001011100000111", -- 5894 FREE #<CONS 0 5895>
 "00000000000000000001011100001000", -- 5895 FREE #<CONS 0 5896>
 "00000000000000000001011100001001", -- 5896 FREE #<CONS 0 5897>
 "00000000000000000001011100001010", -- 5897 FREE #<CONS 0 5898>
 "00000000000000000001011100001011", -- 5898 FREE #<CONS 0 5899>
 "00000000000000000001011100001100", -- 5899 FREE #<CONS 0 5900>
 "00000000000000000001011100001101", -- 5900 FREE #<CONS 0 5901>
 "00000000000000000001011100001110", -- 5901 FREE #<CONS 0 5902>
 "00000000000000000001011100001111", -- 5902 FREE #<CONS 0 5903>
 "00000000000000000001011100010000", -- 5903 FREE #<CONS 0 5904>
 "00000000000000000001011100010001", -- 5904 FREE #<CONS 0 5905>
 "00000000000000000001011100010010", -- 5905 FREE #<CONS 0 5906>
 "00000000000000000001011100010011", -- 5906 FREE #<CONS 0 5907>
 "00000000000000000001011100010100", -- 5907 FREE #<CONS 0 5908>
 "00000000000000000001011100010101", -- 5908 FREE #<CONS 0 5909>
 "00000000000000000001011100010110", -- 5909 FREE #<CONS 0 5910>
 "00000000000000000001011100010111", -- 5910 FREE #<CONS 0 5911>
 "00000000000000000001011100011000", -- 5911 FREE #<CONS 0 5912>
 "00000000000000000001011100011001", -- 5912 FREE #<CONS 0 5913>
 "00000000000000000001011100011010", -- 5913 FREE #<CONS 0 5914>
 "00000000000000000001011100011011", -- 5914 FREE #<CONS 0 5915>
 "00000000000000000001011100011100", -- 5915 FREE #<CONS 0 5916>
 "00000000000000000001011100011101", -- 5916 FREE #<CONS 0 5917>
 "00000000000000000001011100011110", -- 5917 FREE #<CONS 0 5918>
 "00000000000000000001011100011111", -- 5918 FREE #<CONS 0 5919>
 "00000000000000000001011100100000", -- 5919 FREE #<CONS 0 5920>
 "00000000000000000001011100100001", -- 5920 FREE #<CONS 0 5921>
 "00000000000000000001011100100010", -- 5921 FREE #<CONS 0 5922>
 "00000000000000000001011100100011", -- 5922 FREE #<CONS 0 5923>
 "00000000000000000001011100100100", -- 5923 FREE #<CONS 0 5924>
 "00000000000000000001011100100101", -- 5924 FREE #<CONS 0 5925>
 "00000000000000000001011100100110", -- 5925 FREE #<CONS 0 5926>
 "00000000000000000001011100100111", -- 5926 FREE #<CONS 0 5927>
 "00000000000000000001011100101000", -- 5927 FREE #<CONS 0 5928>
 "00000000000000000001011100101001", -- 5928 FREE #<CONS 0 5929>
 "00000000000000000001011100101010", -- 5929 FREE #<CONS 0 5930>
 "00000000000000000001011100101011", -- 5930 FREE #<CONS 0 5931>
 "00000000000000000001011100101100", -- 5931 FREE #<CONS 0 5932>
 "00000000000000000001011100101101", -- 5932 FREE #<CONS 0 5933>
 "00000000000000000001011100101110", -- 5933 FREE #<CONS 0 5934>
 "00000000000000000001011100101111", -- 5934 FREE #<CONS 0 5935>
 "00000000000000000001011100110000", -- 5935 FREE #<CONS 0 5936>
 "00000000000000000001011100110001", -- 5936 FREE #<CONS 0 5937>
 "00000000000000000001011100110010", -- 5937 FREE #<CONS 0 5938>
 "00000000000000000001011100110011", -- 5938 FREE #<CONS 0 5939>
 "00000000000000000001011100110100", -- 5939 FREE #<CONS 0 5940>
 "00000000000000000001011100110101", -- 5940 FREE #<CONS 0 5941>
 "00000000000000000001011100110110", -- 5941 FREE #<CONS 0 5942>
 "00000000000000000001011100110111", -- 5942 FREE #<CONS 0 5943>
 "00000000000000000001011100111000", -- 5943 FREE #<CONS 0 5944>
 "00000000000000000001011100111001", -- 5944 FREE #<CONS 0 5945>
 "00000000000000000001011100111010", -- 5945 FREE #<CONS 0 5946>
 "00000000000000000001011100111011", -- 5946 FREE #<CONS 0 5947>
 "00000000000000000001011100111100", -- 5947 FREE #<CONS 0 5948>
 "00000000000000000001011100111101", -- 5948 FREE #<CONS 0 5949>
 "00000000000000000001011100111110", -- 5949 FREE #<CONS 0 5950>
 "00000000000000000001011100111111", -- 5950 FREE #<CONS 0 5951>
 "00000000000000000001011101000000", -- 5951 FREE #<CONS 0 5952>
 "00000000000000000001011101000001", -- 5952 FREE #<CONS 0 5953>
 "00000000000000000001011101000010", -- 5953 FREE #<CONS 0 5954>
 "00000000000000000001011101000011", -- 5954 FREE #<CONS 0 5955>
 "00000000000000000001011101000100", -- 5955 FREE #<CONS 0 5956>
 "00000000000000000001011101000101", -- 5956 FREE #<CONS 0 5957>
 "00000000000000000001011101000110", -- 5957 FREE #<CONS 0 5958>
 "00000000000000000001011101000111", -- 5958 FREE #<CONS 0 5959>
 "00000000000000000001011101001000", -- 5959 FREE #<CONS 0 5960>
 "00000000000000000001011101001001", -- 5960 FREE #<CONS 0 5961>
 "00000000000000000001011101001010", -- 5961 FREE #<CONS 0 5962>
 "00000000000000000001011101001011", -- 5962 FREE #<CONS 0 5963>
 "00000000000000000001011101001100", -- 5963 FREE #<CONS 0 5964>
 "00000000000000000001011101001101", -- 5964 FREE #<CONS 0 5965>
 "00000000000000000001011101001110", -- 5965 FREE #<CONS 0 5966>
 "00000000000000000001011101001111", -- 5966 FREE #<CONS 0 5967>
 "00000000000000000001011101010000", -- 5967 FREE #<CONS 0 5968>
 "00000000000000000001011101010001", -- 5968 FREE #<CONS 0 5969>
 "00000000000000000001011101010010", -- 5969 FREE #<CONS 0 5970>
 "00000000000000000001011101010011", -- 5970 FREE #<CONS 0 5971>
 "00000000000000000001011101010100", -- 5971 FREE #<CONS 0 5972>
 "00000000000000000001011101010101", -- 5972 FREE #<CONS 0 5973>
 "00000000000000000001011101010110", -- 5973 FREE #<CONS 0 5974>
 "00000000000000000001011101010111", -- 5974 FREE #<CONS 0 5975>
 "00000000000000000001011101011000", -- 5975 FREE #<CONS 0 5976>
 "00000000000000000001011101011001", -- 5976 FREE #<CONS 0 5977>
 "00000000000000000001011101011010", -- 5977 FREE #<CONS 0 5978>
 "00000000000000000001011101011011", -- 5978 FREE #<CONS 0 5979>
 "00000000000000000001011101011100", -- 5979 FREE #<CONS 0 5980>
 "00000000000000000001011101011101", -- 5980 FREE #<CONS 0 5981>
 "00000000000000000001011101011110", -- 5981 FREE #<CONS 0 5982>
 "00000000000000000001011101011111", -- 5982 FREE #<CONS 0 5983>
 "00000000000000000001011101100000", -- 5983 FREE #<CONS 0 5984>
 "00000000000000000001011101100001", -- 5984 FREE #<CONS 0 5985>
 "00000000000000000001011101100010", -- 5985 FREE #<CONS 0 5986>
 "00000000000000000001011101100011", -- 5986 FREE #<CONS 0 5987>
 "00000000000000000001011101100100", -- 5987 FREE #<CONS 0 5988>
 "00000000000000000001011101100101", -- 5988 FREE #<CONS 0 5989>
 "00000000000000000001011101100110", -- 5989 FREE #<CONS 0 5990>
 "00000000000000000001011101100111", -- 5990 FREE #<CONS 0 5991>
 "00000000000000000001011101101000", -- 5991 FREE #<CONS 0 5992>
 "00000000000000000001011101101001", -- 5992 FREE #<CONS 0 5993>
 "00000000000000000001011101101010", -- 5993 FREE #<CONS 0 5994>
 "00000000000000000001011101101011", -- 5994 FREE #<CONS 0 5995>
 "00000000000000000001011101101100", -- 5995 FREE #<CONS 0 5996>
 "00000000000000000001011101101101", -- 5996 FREE #<CONS 0 5997>
 "00000000000000000001011101101110", -- 5997 FREE #<CONS 0 5998>
 "00000000000000000001011101101111", -- 5998 FREE #<CONS 0 5999>
 "00000000000000000001011101110000", -- 5999 FREE #<CONS 0 6000>
 "00000000000000000001011101110001", -- 6000 FREE #<CONS 0 6001>
 "00000000000000000001011101110010", -- 6001 FREE #<CONS 0 6002>
 "00000000000000000001011101110011", -- 6002 FREE #<CONS 0 6003>
 "00000000000000000001011101110100", -- 6003 FREE #<CONS 0 6004>
 "00000000000000000001011101110101", -- 6004 FREE #<CONS 0 6005>
 "00000000000000000001011101110110", -- 6005 FREE #<CONS 0 6006>
 "00000000000000000001011101110111", -- 6006 FREE #<CONS 0 6007>
 "00000000000000000001011101111000", -- 6007 FREE #<CONS 0 6008>
 "00000000000000000001011101111001", -- 6008 FREE #<CONS 0 6009>
 "00000000000000000001011101111010", -- 6009 FREE #<CONS 0 6010>
 "00000000000000000001011101111011", -- 6010 FREE #<CONS 0 6011>
 "00000000000000000001011101111100", -- 6011 FREE #<CONS 0 6012>
 "00000000000000000001011101111101", -- 6012 FREE #<CONS 0 6013>
 "00000000000000000001011101111110", -- 6013 FREE #<CONS 0 6014>
 "00000000000000000001011101111111", -- 6014 FREE #<CONS 0 6015>
 "00000000000000000001011110000000", -- 6015 FREE #<CONS 0 6016>
 "00000000000000000001011110000001", -- 6016 FREE #<CONS 0 6017>
 "00000000000000000001011110000010", -- 6017 FREE #<CONS 0 6018>
 "00000000000000000001011110000011", -- 6018 FREE #<CONS 0 6019>
 "00000000000000000001011110000100", -- 6019 FREE #<CONS 0 6020>
 "00000000000000000001011110000101", -- 6020 FREE #<CONS 0 6021>
 "00000000000000000001011110000110", -- 6021 FREE #<CONS 0 6022>
 "00000000000000000001011110000111", -- 6022 FREE #<CONS 0 6023>
 "00000000000000000001011110001000", -- 6023 FREE #<CONS 0 6024>
 "00000000000000000001011110001001", -- 6024 FREE #<CONS 0 6025>
 "00000000000000000001011110001010", -- 6025 FREE #<CONS 0 6026>
 "00000000000000000001011110001011", -- 6026 FREE #<CONS 0 6027>
 "00000000000000000001011110001100", -- 6027 FREE #<CONS 0 6028>
 "00000000000000000001011110001101", -- 6028 FREE #<CONS 0 6029>
 "00000000000000000001011110001110", -- 6029 FREE #<CONS 0 6030>
 "00000000000000000001011110001111", -- 6030 FREE #<CONS 0 6031>
 "00000000000000000001011110010000", -- 6031 FREE #<CONS 0 6032>
 "00000000000000000001011110010001", -- 6032 FREE #<CONS 0 6033>
 "00000000000000000001011110010010", -- 6033 FREE #<CONS 0 6034>
 "00000000000000000001011110010011", -- 6034 FREE #<CONS 0 6035>
 "00000000000000000001011110010100", -- 6035 FREE #<CONS 0 6036>
 "00000000000000000001011110010101", -- 6036 FREE #<CONS 0 6037>
 "00000000000000000001011110010110", -- 6037 FREE #<CONS 0 6038>
 "00000000000000000001011110010111", -- 6038 FREE #<CONS 0 6039>
 "00000000000000000001011110011000", -- 6039 FREE #<CONS 0 6040>
 "00000000000000000001011110011001", -- 6040 FREE #<CONS 0 6041>
 "00000000000000000001011110011010", -- 6041 FREE #<CONS 0 6042>
 "00000000000000000001011110011011", -- 6042 FREE #<CONS 0 6043>
 "00000000000000000001011110011100", -- 6043 FREE #<CONS 0 6044>
 "00000000000000000001011110011101", -- 6044 FREE #<CONS 0 6045>
 "00000000000000000001011110011110", -- 6045 FREE #<CONS 0 6046>
 "00000000000000000001011110011111", -- 6046 FREE #<CONS 0 6047>
 "00000000000000000001011110100000", -- 6047 FREE #<CONS 0 6048>
 "00000000000000000001011110100001", -- 6048 FREE #<CONS 0 6049>
 "00000000000000000001011110100010", -- 6049 FREE #<CONS 0 6050>
 "00000000000000000001011110100011", -- 6050 FREE #<CONS 0 6051>
 "00000000000000000001011110100100", -- 6051 FREE #<CONS 0 6052>
 "00000000000000000001011110100101", -- 6052 FREE #<CONS 0 6053>
 "00000000000000000001011110100110", -- 6053 FREE #<CONS 0 6054>
 "00000000000000000001011110100111", -- 6054 FREE #<CONS 0 6055>
 "00000000000000000001011110101000", -- 6055 FREE #<CONS 0 6056>
 "00000000000000000001011110101001", -- 6056 FREE #<CONS 0 6057>
 "00000000000000000001011110101010", -- 6057 FREE #<CONS 0 6058>
 "00000000000000000001011110101011", -- 6058 FREE #<CONS 0 6059>
 "00000000000000000001011110101100", -- 6059 FREE #<CONS 0 6060>
 "00000000000000000001011110101101", -- 6060 FREE #<CONS 0 6061>
 "00000000000000000001011110101110", -- 6061 FREE #<CONS 0 6062>
 "00000000000000000001011110101111", -- 6062 FREE #<CONS 0 6063>
 "00000000000000000001011110110000", -- 6063 FREE #<CONS 0 6064>
 "00000000000000000001011110110001", -- 6064 FREE #<CONS 0 6065>
 "00000000000000000001011110110010", -- 6065 FREE #<CONS 0 6066>
 "00000000000000000001011110110011", -- 6066 FREE #<CONS 0 6067>
 "00000000000000000001011110110100", -- 6067 FREE #<CONS 0 6068>
 "00000000000000000001011110110101", -- 6068 FREE #<CONS 0 6069>
 "00000000000000000001011110110110", -- 6069 FREE #<CONS 0 6070>
 "00000000000000000001011110110111", -- 6070 FREE #<CONS 0 6071>
 "00000000000000000001011110111000", -- 6071 FREE #<CONS 0 6072>
 "00000000000000000001011110111001", -- 6072 FREE #<CONS 0 6073>
 "00000000000000000001011110111010", -- 6073 FREE #<CONS 0 6074>
 "00000000000000000001011110111011", -- 6074 FREE #<CONS 0 6075>
 "00000000000000000001011110111100", -- 6075 FREE #<CONS 0 6076>
 "00000000000000000001011110111101", -- 6076 FREE #<CONS 0 6077>
 "00000000000000000001011110111110", -- 6077 FREE #<CONS 0 6078>
 "00000000000000000001011110111111", -- 6078 FREE #<CONS 0 6079>
 "00000000000000000001011111000000", -- 6079 FREE #<CONS 0 6080>
 "00000000000000000001011111000001", -- 6080 FREE #<CONS 0 6081>
 "00000000000000000001011111000010", -- 6081 FREE #<CONS 0 6082>
 "00000000000000000001011111000011", -- 6082 FREE #<CONS 0 6083>
 "00000000000000000001011111000100", -- 6083 FREE #<CONS 0 6084>
 "00000000000000000001011111000101", -- 6084 FREE #<CONS 0 6085>
 "00000000000000000001011111000110", -- 6085 FREE #<CONS 0 6086>
 "00000000000000000001011111000111", -- 6086 FREE #<CONS 0 6087>
 "00000000000000000001011111001000", -- 6087 FREE #<CONS 0 6088>
 "00000000000000000001011111001001", -- 6088 FREE #<CONS 0 6089>
 "00000000000000000001011111001010", -- 6089 FREE #<CONS 0 6090>
 "00000000000000000001011111001011", -- 6090 FREE #<CONS 0 6091>
 "00000000000000000001011111001100", -- 6091 FREE #<CONS 0 6092>
 "00000000000000000001011111001101", -- 6092 FREE #<CONS 0 6093>
 "00000000000000000001011111001110", -- 6093 FREE #<CONS 0 6094>
 "00000000000000000001011111001111", -- 6094 FREE #<CONS 0 6095>
 "00000000000000000001011111010000", -- 6095 FREE #<CONS 0 6096>
 "00000000000000000001011111010001", -- 6096 FREE #<CONS 0 6097>
 "00000000000000000001011111010010", -- 6097 FREE #<CONS 0 6098>
 "00000000000000000001011111010011", -- 6098 FREE #<CONS 0 6099>
 "00000000000000000001011111010100", -- 6099 FREE #<CONS 0 6100>
 "00000000000000000001011111010101", -- 6100 FREE #<CONS 0 6101>
 "00000000000000000001011111010110", -- 6101 FREE #<CONS 0 6102>
 "00000000000000000001011111010111", -- 6102 FREE #<CONS 0 6103>
 "00000000000000000001011111011000", -- 6103 FREE #<CONS 0 6104>
 "00000000000000000001011111011001", -- 6104 FREE #<CONS 0 6105>
 "00000000000000000001011111011010", -- 6105 FREE #<CONS 0 6106>
 "00000000000000000001011111011011", -- 6106 FREE #<CONS 0 6107>
 "00000000000000000001011111011100", -- 6107 FREE #<CONS 0 6108>
 "00000000000000000001011111011101", -- 6108 FREE #<CONS 0 6109>
 "00000000000000000001011111011110", -- 6109 FREE #<CONS 0 6110>
 "00000000000000000001011111011111", -- 6110 FREE #<CONS 0 6111>
 "00000000000000000001011111100000", -- 6111 FREE #<CONS 0 6112>
 "00000000000000000001011111100001", -- 6112 FREE #<CONS 0 6113>
 "00000000000000000001011111100010", -- 6113 FREE #<CONS 0 6114>
 "00000000000000000001011111100011", -- 6114 FREE #<CONS 0 6115>
 "00000000000000000001011111100100", -- 6115 FREE #<CONS 0 6116>
 "00000000000000000001011111100101", -- 6116 FREE #<CONS 0 6117>
 "00000000000000000001011111100110", -- 6117 FREE #<CONS 0 6118>
 "00000000000000000001011111100111", -- 6118 FREE #<CONS 0 6119>
 "00000000000000000001011111101000", -- 6119 FREE #<CONS 0 6120>
 "00000000000000000001011111101001", -- 6120 FREE #<CONS 0 6121>
 "00000000000000000001011111101010", -- 6121 FREE #<CONS 0 6122>
 "00000000000000000001011111101011", -- 6122 FREE #<CONS 0 6123>
 "00000000000000000001011111101100", -- 6123 FREE #<CONS 0 6124>
 "00000000000000000001011111101101", -- 6124 FREE #<CONS 0 6125>
 "00000000000000000001011111101110", -- 6125 FREE #<CONS 0 6126>
 "00000000000000000001011111101111", -- 6126 FREE #<CONS 0 6127>
 "00000000000000000001011111110000", -- 6127 FREE #<CONS 0 6128>
 "00000000000000000001011111110001", -- 6128 FREE #<CONS 0 6129>
 "00000000000000000001011111110010", -- 6129 FREE #<CONS 0 6130>
 "00000000000000000001011111110011", -- 6130 FREE #<CONS 0 6131>
 "00000000000000000001011111110100", -- 6131 FREE #<CONS 0 6132>
 "00000000000000000001011111110101", -- 6132 FREE #<CONS 0 6133>
 "00000000000000000001011111110110", -- 6133 FREE #<CONS 0 6134>
 "00000000000000000001011111110111", -- 6134 FREE #<CONS 0 6135>
 "00000000000000000001011111111000", -- 6135 FREE #<CONS 0 6136>
 "00000000000000000001011111111001", -- 6136 FREE #<CONS 0 6137>
 "00000000000000000001011111111010", -- 6137 FREE #<CONS 0 6138>
 "00000000000000000001011111111011", -- 6138 FREE #<CONS 0 6139>
 "00000000000000000001011111111100", -- 6139 FREE #<CONS 0 6140>
 "00000000000000000001011111111101", -- 6140 FREE #<CONS 0 6141>
 "00000000000000000001011111111110", -- 6141 FREE #<CONS 0 6142>
 "00000000000000000001011111111111", -- 6142 FREE #<CONS 0 6143>
 "00000000000000000001100000000000", -- 6143 FREE #<CONS 0 6144>
 "00000000000000000001100000000001", -- 6144 FREE #<CONS 0 6145>
 "00000000000000000001100000000010", -- 6145 FREE #<CONS 0 6146>
 "00000000000000000001100000000011", -- 6146 FREE #<CONS 0 6147>
 "00000000000000000001100000000100", -- 6147 FREE #<CONS 0 6148>
 "00000000000000000001100000000101", -- 6148 FREE #<CONS 0 6149>
 "00000000000000000001100000000110", -- 6149 FREE #<CONS 0 6150>
 "00000000000000000001100000000111", -- 6150 FREE #<CONS 0 6151>
 "00000000000000000001100000001000", -- 6151 FREE #<CONS 0 6152>
 "00000000000000000001100000001001", -- 6152 FREE #<CONS 0 6153>
 "00000000000000000001100000001010", -- 6153 FREE #<CONS 0 6154>
 "00000000000000000001100000001011", -- 6154 FREE #<CONS 0 6155>
 "00000000000000000001100000001100", -- 6155 FREE #<CONS 0 6156>
 "00000000000000000001100000001101", -- 6156 FREE #<CONS 0 6157>
 "00000000000000000001100000001110", -- 6157 FREE #<CONS 0 6158>
 "00000000000000000001100000001111", -- 6158 FREE #<CONS 0 6159>
 "00000000000000000001100000010000", -- 6159 FREE #<CONS 0 6160>
 "00000000000000000001100000010001", -- 6160 FREE #<CONS 0 6161>
 "00000000000000000001100000010010", -- 6161 FREE #<CONS 0 6162>
 "00000000000000000001100000010011", -- 6162 FREE #<CONS 0 6163>
 "00000000000000000001100000010100", -- 6163 FREE #<CONS 0 6164>
 "00000000000000000001100000010101", -- 6164 FREE #<CONS 0 6165>
 "00000000000000000001100000010110", -- 6165 FREE #<CONS 0 6166>
 "00000000000000000001100000010111", -- 6166 FREE #<CONS 0 6167>
 "00000000000000000001100000011000", -- 6167 FREE #<CONS 0 6168>
 "00000000000000000001100000011001", -- 6168 FREE #<CONS 0 6169>
 "00000000000000000001100000011010", -- 6169 FREE #<CONS 0 6170>
 "00000000000000000001100000011011", -- 6170 FREE #<CONS 0 6171>
 "00000000000000000001100000011100", -- 6171 FREE #<CONS 0 6172>
 "00000000000000000001100000011101", -- 6172 FREE #<CONS 0 6173>
 "00000000000000000001100000011110", -- 6173 FREE #<CONS 0 6174>
 "00000000000000000001100000011111", -- 6174 FREE #<CONS 0 6175>
 "00000000000000000001100000100000", -- 6175 FREE #<CONS 0 6176>
 "00000000000000000001100000100001", -- 6176 FREE #<CONS 0 6177>
 "00000000000000000001100000100010", -- 6177 FREE #<CONS 0 6178>
 "00000000000000000001100000100011", -- 6178 FREE #<CONS 0 6179>
 "00000000000000000001100000100100", -- 6179 FREE #<CONS 0 6180>
 "00000000000000000001100000100101", -- 6180 FREE #<CONS 0 6181>
 "00000000000000000001100000100110", -- 6181 FREE #<CONS 0 6182>
 "00000000000000000001100000100111", -- 6182 FREE #<CONS 0 6183>
 "00000000000000000001100000101000", -- 6183 FREE #<CONS 0 6184>
 "00000000000000000001100000101001", -- 6184 FREE #<CONS 0 6185>
 "00000000000000000001100000101010", -- 6185 FREE #<CONS 0 6186>
 "00000000000000000001100000101011", -- 6186 FREE #<CONS 0 6187>
 "00000000000000000001100000101100", -- 6187 FREE #<CONS 0 6188>
 "00000000000000000001100000101101", -- 6188 FREE #<CONS 0 6189>
 "00000000000000000001100000101110", -- 6189 FREE #<CONS 0 6190>
 "00000000000000000001100000101111", -- 6190 FREE #<CONS 0 6191>
 "00000000000000000001100000110000", -- 6191 FREE #<CONS 0 6192>
 "00000000000000000001100000110001", -- 6192 FREE #<CONS 0 6193>
 "00000000000000000001100000110010", -- 6193 FREE #<CONS 0 6194>
 "00000000000000000001100000110011", -- 6194 FREE #<CONS 0 6195>
 "00000000000000000001100000110100", -- 6195 FREE #<CONS 0 6196>
 "00000000000000000001100000110101", -- 6196 FREE #<CONS 0 6197>
 "00000000000000000001100000110110", -- 6197 FREE #<CONS 0 6198>
 "00000000000000000001100000110111", -- 6198 FREE #<CONS 0 6199>
 "00000000000000000001100000111000", -- 6199 FREE #<CONS 0 6200>
 "00000000000000000001100000111001", -- 6200 FREE #<CONS 0 6201>
 "00000000000000000001100000111010", -- 6201 FREE #<CONS 0 6202>
 "00000000000000000001100000111011", -- 6202 FREE #<CONS 0 6203>
 "00000000000000000001100000111100", -- 6203 FREE #<CONS 0 6204>
 "00000000000000000001100000111101", -- 6204 FREE #<CONS 0 6205>
 "00000000000000000001100000111110", -- 6205 FREE #<CONS 0 6206>
 "00000000000000000001100000111111", -- 6206 FREE #<CONS 0 6207>
 "00000000000000000001100001000000", -- 6207 FREE #<CONS 0 6208>
 "00000000000000000001100001000001", -- 6208 FREE #<CONS 0 6209>
 "00000000000000000001100001000010", -- 6209 FREE #<CONS 0 6210>
 "00000000000000000001100001000011", -- 6210 FREE #<CONS 0 6211>
 "00000000000000000001100001000100", -- 6211 FREE #<CONS 0 6212>
 "00000000000000000001100001000101", -- 6212 FREE #<CONS 0 6213>
 "00000000000000000001100001000110", -- 6213 FREE #<CONS 0 6214>
 "00000000000000000001100001000111", -- 6214 FREE #<CONS 0 6215>
 "00000000000000000001100001001000", -- 6215 FREE #<CONS 0 6216>
 "00000000000000000001100001001001", -- 6216 FREE #<CONS 0 6217>
 "00000000000000000001100001001010", -- 6217 FREE #<CONS 0 6218>
 "00000000000000000001100001001011", -- 6218 FREE #<CONS 0 6219>
 "00000000000000000001100001001100", -- 6219 FREE #<CONS 0 6220>
 "00000000000000000001100001001101", -- 6220 FREE #<CONS 0 6221>
 "00000000000000000001100001001110", -- 6221 FREE #<CONS 0 6222>
 "00000000000000000001100001001111", -- 6222 FREE #<CONS 0 6223>
 "00000000000000000001100001010000", -- 6223 FREE #<CONS 0 6224>
 "00000000000000000001100001010001", -- 6224 FREE #<CONS 0 6225>
 "00000000000000000001100001010010", -- 6225 FREE #<CONS 0 6226>
 "00000000000000000001100001010011", -- 6226 FREE #<CONS 0 6227>
 "00000000000000000001100001010100", -- 6227 FREE #<CONS 0 6228>
 "00000000000000000001100001010101", -- 6228 FREE #<CONS 0 6229>
 "00000000000000000001100001010110", -- 6229 FREE #<CONS 0 6230>
 "00000000000000000001100001010111", -- 6230 FREE #<CONS 0 6231>
 "00000000000000000001100001011000", -- 6231 FREE #<CONS 0 6232>
 "00000000000000000001100001011001", -- 6232 FREE #<CONS 0 6233>
 "00000000000000000001100001011010", -- 6233 FREE #<CONS 0 6234>
 "00000000000000000001100001011011", -- 6234 FREE #<CONS 0 6235>
 "00000000000000000001100001011100", -- 6235 FREE #<CONS 0 6236>
 "00000000000000000001100001011101", -- 6236 FREE #<CONS 0 6237>
 "00000000000000000001100001011110", -- 6237 FREE #<CONS 0 6238>
 "00000000000000000001100001011111", -- 6238 FREE #<CONS 0 6239>
 "00000000000000000001100001100000", -- 6239 FREE #<CONS 0 6240>
 "00000000000000000001100001100001", -- 6240 FREE #<CONS 0 6241>
 "00000000000000000001100001100010", -- 6241 FREE #<CONS 0 6242>
 "00000000000000000001100001100011", -- 6242 FREE #<CONS 0 6243>
 "00000000000000000001100001100100", -- 6243 FREE #<CONS 0 6244>
 "00000000000000000001100001100101", -- 6244 FREE #<CONS 0 6245>
 "00000000000000000001100001100110", -- 6245 FREE #<CONS 0 6246>
 "00000000000000000001100001100111", -- 6246 FREE #<CONS 0 6247>
 "00000000000000000001100001101000", -- 6247 FREE #<CONS 0 6248>
 "00000000000000000001100001101001", -- 6248 FREE #<CONS 0 6249>
 "00000000000000000001100001101010", -- 6249 FREE #<CONS 0 6250>
 "00000000000000000001100001101011", -- 6250 FREE #<CONS 0 6251>
 "00000000000000000001100001101100", -- 6251 FREE #<CONS 0 6252>
 "00000000000000000001100001101101", -- 6252 FREE #<CONS 0 6253>
 "00000000000000000001100001101110", -- 6253 FREE #<CONS 0 6254>
 "00000000000000000001100001101111", -- 6254 FREE #<CONS 0 6255>
 "00000000000000000001100001110000", -- 6255 FREE #<CONS 0 6256>
 "00000000000000000001100001110001", -- 6256 FREE #<CONS 0 6257>
 "00000000000000000001100001110010", -- 6257 FREE #<CONS 0 6258>
 "00000000000000000001100001110011", -- 6258 FREE #<CONS 0 6259>
 "00000000000000000001100001110100", -- 6259 FREE #<CONS 0 6260>
 "00000000000000000001100001110101", -- 6260 FREE #<CONS 0 6261>
 "00000000000000000001100001110110", -- 6261 FREE #<CONS 0 6262>
 "00000000000000000001100001110111", -- 6262 FREE #<CONS 0 6263>
 "00000000000000000001100001111000", -- 6263 FREE #<CONS 0 6264>
 "00000000000000000001100001111001", -- 6264 FREE #<CONS 0 6265>
 "00000000000000000001100001111010", -- 6265 FREE #<CONS 0 6266>
 "00000000000000000001100001111011", -- 6266 FREE #<CONS 0 6267>
 "00000000000000000001100001111100", -- 6267 FREE #<CONS 0 6268>
 "00000000000000000001100001111101", -- 6268 FREE #<CONS 0 6269>
 "00000000000000000001100001111110", -- 6269 FREE #<CONS 0 6270>
 "00000000000000000001100001111111", -- 6270 FREE #<CONS 0 6271>
 "00000000000000000001100010000000", -- 6271 FREE #<CONS 0 6272>
 "00000000000000000001100010000001", -- 6272 FREE #<CONS 0 6273>
 "00000000000000000001100010000010", -- 6273 FREE #<CONS 0 6274>
 "00000000000000000001100010000011", -- 6274 FREE #<CONS 0 6275>
 "00000000000000000001100010000100", -- 6275 FREE #<CONS 0 6276>
 "00000000000000000001100010000101", -- 6276 FREE #<CONS 0 6277>
 "00000000000000000001100010000110", -- 6277 FREE #<CONS 0 6278>
 "00000000000000000001100010000111", -- 6278 FREE #<CONS 0 6279>
 "00000000000000000001100010001000", -- 6279 FREE #<CONS 0 6280>
 "00000000000000000001100010001001", -- 6280 FREE #<CONS 0 6281>
 "00000000000000000001100010001010", -- 6281 FREE #<CONS 0 6282>
 "00000000000000000001100010001011", -- 6282 FREE #<CONS 0 6283>
 "00000000000000000001100010001100", -- 6283 FREE #<CONS 0 6284>
 "00000000000000000001100010001101", -- 6284 FREE #<CONS 0 6285>
 "00000000000000000001100010001110", -- 6285 FREE #<CONS 0 6286>
 "00000000000000000001100010001111", -- 6286 FREE #<CONS 0 6287>
 "00000000000000000001100010010000", -- 6287 FREE #<CONS 0 6288>
 "00000000000000000001100010010001", -- 6288 FREE #<CONS 0 6289>
 "00000000000000000001100010010010", -- 6289 FREE #<CONS 0 6290>
 "00000000000000000001100010010011", -- 6290 FREE #<CONS 0 6291>
 "00000000000000000001100010010100", -- 6291 FREE #<CONS 0 6292>
 "00000000000000000001100010010101", -- 6292 FREE #<CONS 0 6293>
 "00000000000000000001100010010110", -- 6293 FREE #<CONS 0 6294>
 "00000000000000000001100010010111", -- 6294 FREE #<CONS 0 6295>
 "00000000000000000001100010011000", -- 6295 FREE #<CONS 0 6296>
 "00000000000000000001100010011001", -- 6296 FREE #<CONS 0 6297>
 "00000000000000000001100010011010", -- 6297 FREE #<CONS 0 6298>
 "00000000000000000001100010011011", -- 6298 FREE #<CONS 0 6299>
 "00000000000000000001100010011100", -- 6299 FREE #<CONS 0 6300>
 "00000000000000000001100010011101", -- 6300 FREE #<CONS 0 6301>
 "00000000000000000001100010011110", -- 6301 FREE #<CONS 0 6302>
 "00000000000000000001100010011111", -- 6302 FREE #<CONS 0 6303>
 "00000000000000000001100010100000", -- 6303 FREE #<CONS 0 6304>
 "00000000000000000001100010100001", -- 6304 FREE #<CONS 0 6305>
 "00000000000000000001100010100010", -- 6305 FREE #<CONS 0 6306>
 "00000000000000000001100010100011", -- 6306 FREE #<CONS 0 6307>
 "00000000000000000001100010100100", -- 6307 FREE #<CONS 0 6308>
 "00000000000000000001100010100101", -- 6308 FREE #<CONS 0 6309>
 "00000000000000000001100010100110", -- 6309 FREE #<CONS 0 6310>
 "00000000000000000001100010100111", -- 6310 FREE #<CONS 0 6311>
 "00000000000000000001100010101000", -- 6311 FREE #<CONS 0 6312>
 "00000000000000000001100010101001", -- 6312 FREE #<CONS 0 6313>
 "00000000000000000001100010101010", -- 6313 FREE #<CONS 0 6314>
 "00000000000000000001100010101011", -- 6314 FREE #<CONS 0 6315>
 "00000000000000000001100010101100", -- 6315 FREE #<CONS 0 6316>
 "00000000000000000001100010101101", -- 6316 FREE #<CONS 0 6317>
 "00000000000000000001100010101110", -- 6317 FREE #<CONS 0 6318>
 "00000000000000000001100010101111", -- 6318 FREE #<CONS 0 6319>
 "00000000000000000001100010110000", -- 6319 FREE #<CONS 0 6320>
 "00000000000000000001100010110001", -- 6320 FREE #<CONS 0 6321>
 "00000000000000000001100010110010", -- 6321 FREE #<CONS 0 6322>
 "00000000000000000001100010110011", -- 6322 FREE #<CONS 0 6323>
 "00000000000000000001100010110100", -- 6323 FREE #<CONS 0 6324>
 "00000000000000000001100010110101", -- 6324 FREE #<CONS 0 6325>
 "00000000000000000001100010110110", -- 6325 FREE #<CONS 0 6326>
 "00000000000000000001100010110111", -- 6326 FREE #<CONS 0 6327>
 "00000000000000000001100010111000", -- 6327 FREE #<CONS 0 6328>
 "00000000000000000001100010111001", -- 6328 FREE #<CONS 0 6329>
 "00000000000000000001100010111010", -- 6329 FREE #<CONS 0 6330>
 "00000000000000000001100010111011", -- 6330 FREE #<CONS 0 6331>
 "00000000000000000001100010111100", -- 6331 FREE #<CONS 0 6332>
 "00000000000000000001100010111101", -- 6332 FREE #<CONS 0 6333>
 "00000000000000000001100010111110", -- 6333 FREE #<CONS 0 6334>
 "00000000000000000001100010111111", -- 6334 FREE #<CONS 0 6335>
 "00000000000000000001100011000000", -- 6335 FREE #<CONS 0 6336>
 "00000000000000000001100011000001", -- 6336 FREE #<CONS 0 6337>
 "00000000000000000001100011000010", -- 6337 FREE #<CONS 0 6338>
 "00000000000000000001100011000011", -- 6338 FREE #<CONS 0 6339>
 "00000000000000000001100011000100", -- 6339 FREE #<CONS 0 6340>
 "00000000000000000001100011000101", -- 6340 FREE #<CONS 0 6341>
 "00000000000000000001100011000110", -- 6341 FREE #<CONS 0 6342>
 "00000000000000000001100011000111", -- 6342 FREE #<CONS 0 6343>
 "00000000000000000001100011001000", -- 6343 FREE #<CONS 0 6344>
 "00000000000000000001100011001001", -- 6344 FREE #<CONS 0 6345>
 "00000000000000000001100011001010", -- 6345 FREE #<CONS 0 6346>
 "00000000000000000001100011001011", -- 6346 FREE #<CONS 0 6347>
 "00000000000000000001100011001100", -- 6347 FREE #<CONS 0 6348>
 "00000000000000000001100011001101", -- 6348 FREE #<CONS 0 6349>
 "00000000000000000001100011001110", -- 6349 FREE #<CONS 0 6350>
 "00000000000000000001100011001111", -- 6350 FREE #<CONS 0 6351>
 "00000000000000000001100011010000", -- 6351 FREE #<CONS 0 6352>
 "00000000000000000001100011010001", -- 6352 FREE #<CONS 0 6353>
 "00000000000000000001100011010010", -- 6353 FREE #<CONS 0 6354>
 "00000000000000000001100011010011", -- 6354 FREE #<CONS 0 6355>
 "00000000000000000001100011010100", -- 6355 FREE #<CONS 0 6356>
 "00000000000000000001100011010101", -- 6356 FREE #<CONS 0 6357>
 "00000000000000000001100011010110", -- 6357 FREE #<CONS 0 6358>
 "00000000000000000001100011010111", -- 6358 FREE #<CONS 0 6359>
 "00000000000000000001100011011000", -- 6359 FREE #<CONS 0 6360>
 "00000000000000000001100011011001", -- 6360 FREE #<CONS 0 6361>
 "00000000000000000001100011011010", -- 6361 FREE #<CONS 0 6362>
 "00000000000000000001100011011011", -- 6362 FREE #<CONS 0 6363>
 "00000000000000000001100011011100", -- 6363 FREE #<CONS 0 6364>
 "00000000000000000001100011011101", -- 6364 FREE #<CONS 0 6365>
 "00000000000000000001100011011110", -- 6365 FREE #<CONS 0 6366>
 "00000000000000000001100011011111", -- 6366 FREE #<CONS 0 6367>
 "00000000000000000001100011100000", -- 6367 FREE #<CONS 0 6368>
 "00000000000000000001100011100001", -- 6368 FREE #<CONS 0 6369>
 "00000000000000000001100011100010", -- 6369 FREE #<CONS 0 6370>
 "00000000000000000001100011100011", -- 6370 FREE #<CONS 0 6371>
 "00000000000000000001100011100100", -- 6371 FREE #<CONS 0 6372>
 "00000000000000000001100011100101", -- 6372 FREE #<CONS 0 6373>
 "00000000000000000001100011100110", -- 6373 FREE #<CONS 0 6374>
 "00000000000000000001100011100111", -- 6374 FREE #<CONS 0 6375>
 "00000000000000000001100011101000", -- 6375 FREE #<CONS 0 6376>
 "00000000000000000001100011101001", -- 6376 FREE #<CONS 0 6377>
 "00000000000000000001100011101010", -- 6377 FREE #<CONS 0 6378>
 "00000000000000000001100011101011", -- 6378 FREE #<CONS 0 6379>
 "00000000000000000001100011101100", -- 6379 FREE #<CONS 0 6380>
 "00000000000000000001100011101101", -- 6380 FREE #<CONS 0 6381>
 "00000000000000000001100011101110", -- 6381 FREE #<CONS 0 6382>
 "00000000000000000001100011101111", -- 6382 FREE #<CONS 0 6383>
 "00000000000000000001100011110000", -- 6383 FREE #<CONS 0 6384>
 "00000000000000000001100011110001", -- 6384 FREE #<CONS 0 6385>
 "00000000000000000001100011110010", -- 6385 FREE #<CONS 0 6386>
 "00000000000000000001100011110011", -- 6386 FREE #<CONS 0 6387>
 "00000000000000000001100011110100", -- 6387 FREE #<CONS 0 6388>
 "00000000000000000001100011110101", -- 6388 FREE #<CONS 0 6389>
 "00000000000000000001100011110110", -- 6389 FREE #<CONS 0 6390>
 "00000000000000000001100011110111", -- 6390 FREE #<CONS 0 6391>
 "00000000000000000001100011111000", -- 6391 FREE #<CONS 0 6392>
 "00000000000000000001100011111001", -- 6392 FREE #<CONS 0 6393>
 "00000000000000000001100011111010", -- 6393 FREE #<CONS 0 6394>
 "00000000000000000001100011111011", -- 6394 FREE #<CONS 0 6395>
 "00000000000000000001100011111100", -- 6395 FREE #<CONS 0 6396>
 "00000000000000000001100011111101", -- 6396 FREE #<CONS 0 6397>
 "00000000000000000001100011111110", -- 6397 FREE #<CONS 0 6398>
 "00000000000000000001100011111111", -- 6398 FREE #<CONS 0 6399>
 "00000000000000000001100100000000", -- 6399 FREE #<CONS 0 6400>
 "00000000000000000001100100000001", -- 6400 FREE #<CONS 0 6401>
 "00000000000000000001100100000010", -- 6401 FREE #<CONS 0 6402>
 "00000000000000000001100100000011", -- 6402 FREE #<CONS 0 6403>
 "00000000000000000001100100000100", -- 6403 FREE #<CONS 0 6404>
 "00000000000000000001100100000101", -- 6404 FREE #<CONS 0 6405>
 "00000000000000000001100100000110", -- 6405 FREE #<CONS 0 6406>
 "00000000000000000001100100000111", -- 6406 FREE #<CONS 0 6407>
 "00000000000000000001100100001000", -- 6407 FREE #<CONS 0 6408>
 "00000000000000000001100100001001", -- 6408 FREE #<CONS 0 6409>
 "00000000000000000001100100001010", -- 6409 FREE #<CONS 0 6410>
 "00000000000000000001100100001011", -- 6410 FREE #<CONS 0 6411>
 "00000000000000000001100100001100", -- 6411 FREE #<CONS 0 6412>
 "00000000000000000001100100001101", -- 6412 FREE #<CONS 0 6413>
 "00000000000000000001100100001110", -- 6413 FREE #<CONS 0 6414>
 "00000000000000000001100100001111", -- 6414 FREE #<CONS 0 6415>
 "00000000000000000001100100010000", -- 6415 FREE #<CONS 0 6416>
 "00000000000000000001100100010001", -- 6416 FREE #<CONS 0 6417>
 "00000000000000000001100100010010", -- 6417 FREE #<CONS 0 6418>
 "00000000000000000001100100010011", -- 6418 FREE #<CONS 0 6419>
 "00000000000000000001100100010100", -- 6419 FREE #<CONS 0 6420>
 "00000000000000000001100100010101", -- 6420 FREE #<CONS 0 6421>
 "00000000000000000001100100010110", -- 6421 FREE #<CONS 0 6422>
 "00000000000000000001100100010111", -- 6422 FREE #<CONS 0 6423>
 "00000000000000000001100100011000", -- 6423 FREE #<CONS 0 6424>
 "00000000000000000001100100011001", -- 6424 FREE #<CONS 0 6425>
 "00000000000000000001100100011010", -- 6425 FREE #<CONS 0 6426>
 "00000000000000000001100100011011", -- 6426 FREE #<CONS 0 6427>
 "00000000000000000001100100011100", -- 6427 FREE #<CONS 0 6428>
 "00000000000000000001100100011101", -- 6428 FREE #<CONS 0 6429>
 "00000000000000000001100100011110", -- 6429 FREE #<CONS 0 6430>
 "00000000000000000001100100011111", -- 6430 FREE #<CONS 0 6431>
 "00000000000000000001100100100000", -- 6431 FREE #<CONS 0 6432>
 "00000000000000000001100100100001", -- 6432 FREE #<CONS 0 6433>
 "00000000000000000001100100100010", -- 6433 FREE #<CONS 0 6434>
 "00000000000000000001100100100011", -- 6434 FREE #<CONS 0 6435>
 "00000000000000000001100100100100", -- 6435 FREE #<CONS 0 6436>
 "00000000000000000001100100100101", -- 6436 FREE #<CONS 0 6437>
 "00000000000000000001100100100110", -- 6437 FREE #<CONS 0 6438>
 "00000000000000000001100100100111", -- 6438 FREE #<CONS 0 6439>
 "00000000000000000001100100101000", -- 6439 FREE #<CONS 0 6440>
 "00000000000000000001100100101001", -- 6440 FREE #<CONS 0 6441>
 "00000000000000000001100100101010", -- 6441 FREE #<CONS 0 6442>
 "00000000000000000001100100101011", -- 6442 FREE #<CONS 0 6443>
 "00000000000000000001100100101100", -- 6443 FREE #<CONS 0 6444>
 "00000000000000000001100100101101", -- 6444 FREE #<CONS 0 6445>
 "00000000000000000001100100101110", -- 6445 FREE #<CONS 0 6446>
 "00000000000000000001100100101111", -- 6446 FREE #<CONS 0 6447>
 "00000000000000000001100100110000", -- 6447 FREE #<CONS 0 6448>
 "00000000000000000001100100110001", -- 6448 FREE #<CONS 0 6449>
 "00000000000000000001100100110010", -- 6449 FREE #<CONS 0 6450>
 "00000000000000000001100100110011", -- 6450 FREE #<CONS 0 6451>
 "00000000000000000001100100110100", -- 6451 FREE #<CONS 0 6452>
 "00000000000000000001100100110101", -- 6452 FREE #<CONS 0 6453>
 "00000000000000000001100100110110", -- 6453 FREE #<CONS 0 6454>
 "00000000000000000001100100110111", -- 6454 FREE #<CONS 0 6455>
 "00000000000000000001100100111000", -- 6455 FREE #<CONS 0 6456>
 "00000000000000000001100100111001", -- 6456 FREE #<CONS 0 6457>
 "00000000000000000001100100111010", -- 6457 FREE #<CONS 0 6458>
 "00000000000000000001100100111011", -- 6458 FREE #<CONS 0 6459>
 "00000000000000000001100100111100", -- 6459 FREE #<CONS 0 6460>
 "00000000000000000001100100111101", -- 6460 FREE #<CONS 0 6461>
 "00000000000000000001100100111110", -- 6461 FREE #<CONS 0 6462>
 "00000000000000000001100100111111", -- 6462 FREE #<CONS 0 6463>
 "00000000000000000001100101000000", -- 6463 FREE #<CONS 0 6464>
 "00000000000000000001100101000001", -- 6464 FREE #<CONS 0 6465>
 "00000000000000000001100101000010", -- 6465 FREE #<CONS 0 6466>
 "00000000000000000001100101000011", -- 6466 FREE #<CONS 0 6467>
 "00000000000000000001100101000100", -- 6467 FREE #<CONS 0 6468>
 "00000000000000000001100101000101", -- 6468 FREE #<CONS 0 6469>
 "00000000000000000001100101000110", -- 6469 FREE #<CONS 0 6470>
 "00000000000000000001100101000111", -- 6470 FREE #<CONS 0 6471>
 "00000000000000000001100101001000", -- 6471 FREE #<CONS 0 6472>
 "00000000000000000001100101001001", -- 6472 FREE #<CONS 0 6473>
 "00000000000000000001100101001010", -- 6473 FREE #<CONS 0 6474>
 "00000000000000000001100101001011", -- 6474 FREE #<CONS 0 6475>
 "00000000000000000001100101001100", -- 6475 FREE #<CONS 0 6476>
 "00000000000000000001100101001101", -- 6476 FREE #<CONS 0 6477>
 "00000000000000000001100101001110", -- 6477 FREE #<CONS 0 6478>
 "00000000000000000001100101001111", -- 6478 FREE #<CONS 0 6479>
 "00000000000000000001100101010000", -- 6479 FREE #<CONS 0 6480>
 "00000000000000000001100101010001", -- 6480 FREE #<CONS 0 6481>
 "00000000000000000001100101010010", -- 6481 FREE #<CONS 0 6482>
 "00000000000000000001100101010011", -- 6482 FREE #<CONS 0 6483>
 "00000000000000000001100101010100", -- 6483 FREE #<CONS 0 6484>
 "00000000000000000001100101010101", -- 6484 FREE #<CONS 0 6485>
 "00000000000000000001100101010110", -- 6485 FREE #<CONS 0 6486>
 "00000000000000000001100101010111", -- 6486 FREE #<CONS 0 6487>
 "00000000000000000001100101011000", -- 6487 FREE #<CONS 0 6488>
 "00000000000000000001100101011001", -- 6488 FREE #<CONS 0 6489>
 "00000000000000000001100101011010", -- 6489 FREE #<CONS 0 6490>
 "00000000000000000001100101011011", -- 6490 FREE #<CONS 0 6491>
 "00000000000000000001100101011100", -- 6491 FREE #<CONS 0 6492>
 "00000000000000000001100101011101", -- 6492 FREE #<CONS 0 6493>
 "00000000000000000001100101011110", -- 6493 FREE #<CONS 0 6494>
 "00000000000000000001100101011111", -- 6494 FREE #<CONS 0 6495>
 "00000000000000000001100101100000", -- 6495 FREE #<CONS 0 6496>
 "00000000000000000001100101100001", -- 6496 FREE #<CONS 0 6497>
 "00000000000000000001100101100010", -- 6497 FREE #<CONS 0 6498>
 "00000000000000000001100101100011", -- 6498 FREE #<CONS 0 6499>
 "00000000000000000001100101100100", -- 6499 FREE #<CONS 0 6500>
 "00000000000000000001100101100101", -- 6500 FREE #<CONS 0 6501>
 "00000000000000000001100101100110", -- 6501 FREE #<CONS 0 6502>
 "00000000000000000001100101100111", -- 6502 FREE #<CONS 0 6503>
 "00000000000000000001100101101000", -- 6503 FREE #<CONS 0 6504>
 "00000000000000000001100101101001", -- 6504 FREE #<CONS 0 6505>
 "00000000000000000001100101101010", -- 6505 FREE #<CONS 0 6506>
 "00000000000000000001100101101011", -- 6506 FREE #<CONS 0 6507>
 "00000000000000000001100101101100", -- 6507 FREE #<CONS 0 6508>
 "00000000000000000001100101101101", -- 6508 FREE #<CONS 0 6509>
 "00000000000000000001100101101110", -- 6509 FREE #<CONS 0 6510>
 "00000000000000000001100101101111", -- 6510 FREE #<CONS 0 6511>
 "00000000000000000001100101110000", -- 6511 FREE #<CONS 0 6512>
 "00000000000000000001100101110001", -- 6512 FREE #<CONS 0 6513>
 "00000000000000000001100101110010", -- 6513 FREE #<CONS 0 6514>
 "00000000000000000001100101110011", -- 6514 FREE #<CONS 0 6515>
 "00000000000000000001100101110100", -- 6515 FREE #<CONS 0 6516>
 "00000000000000000001100101110101", -- 6516 FREE #<CONS 0 6517>
 "00000000000000000001100101110110", -- 6517 FREE #<CONS 0 6518>
 "00000000000000000001100101110111", -- 6518 FREE #<CONS 0 6519>
 "00000000000000000001100101111000", -- 6519 FREE #<CONS 0 6520>
 "00000000000000000001100101111001", -- 6520 FREE #<CONS 0 6521>
 "00000000000000000001100101111010", -- 6521 FREE #<CONS 0 6522>
 "00000000000000000001100101111011", -- 6522 FREE #<CONS 0 6523>
 "00000000000000000001100101111100", -- 6523 FREE #<CONS 0 6524>
 "00000000000000000001100101111101", -- 6524 FREE #<CONS 0 6525>
 "00000000000000000001100101111110", -- 6525 FREE #<CONS 0 6526>
 "00000000000000000001100101111111", -- 6526 FREE #<CONS 0 6527>
 "00000000000000000001100110000000", -- 6527 FREE #<CONS 0 6528>
 "00000000000000000001100110000001", -- 6528 FREE #<CONS 0 6529>
 "00000000000000000001100110000010", -- 6529 FREE #<CONS 0 6530>
 "00000000000000000001100110000011", -- 6530 FREE #<CONS 0 6531>
 "00000000000000000001100110000100", -- 6531 FREE #<CONS 0 6532>
 "00000000000000000001100110000101", -- 6532 FREE #<CONS 0 6533>
 "00000000000000000001100110000110", -- 6533 FREE #<CONS 0 6534>
 "00000000000000000001100110000111", -- 6534 FREE #<CONS 0 6535>
 "00000000000000000001100110001000", -- 6535 FREE #<CONS 0 6536>
 "00000000000000000001100110001001", -- 6536 FREE #<CONS 0 6537>
 "00000000000000000001100110001010", -- 6537 FREE #<CONS 0 6538>
 "00000000000000000001100110001011", -- 6538 FREE #<CONS 0 6539>
 "00000000000000000001100110001100", -- 6539 FREE #<CONS 0 6540>
 "00000000000000000001100110001101", -- 6540 FREE #<CONS 0 6541>
 "00000000000000000001100110001110", -- 6541 FREE #<CONS 0 6542>
 "00000000000000000001100110001111", -- 6542 FREE #<CONS 0 6543>
 "00000000000000000001100110010000", -- 6543 FREE #<CONS 0 6544>
 "00000000000000000001100110010001", -- 6544 FREE #<CONS 0 6545>
 "00000000000000000001100110010010", -- 6545 FREE #<CONS 0 6546>
 "00000000000000000001100110010011", -- 6546 FREE #<CONS 0 6547>
 "00000000000000000001100110010100", -- 6547 FREE #<CONS 0 6548>
 "00000000000000000001100110010101", -- 6548 FREE #<CONS 0 6549>
 "00000000000000000001100110010110", -- 6549 FREE #<CONS 0 6550>
 "00000000000000000001100110010111", -- 6550 FREE #<CONS 0 6551>
 "00000000000000000001100110011000", -- 6551 FREE #<CONS 0 6552>
 "00000000000000000001100110011001", -- 6552 FREE #<CONS 0 6553>
 "00000000000000000001100110011010", -- 6553 FREE #<CONS 0 6554>
 "00000000000000000001100110011011", -- 6554 FREE #<CONS 0 6555>
 "00000000000000000001100110011100", -- 6555 FREE #<CONS 0 6556>
 "00000000000000000001100110011101", -- 6556 FREE #<CONS 0 6557>
 "00000000000000000001100110011110", -- 6557 FREE #<CONS 0 6558>
 "00000000000000000001100110011111", -- 6558 FREE #<CONS 0 6559>
 "00000000000000000001100110100000", -- 6559 FREE #<CONS 0 6560>
 "00000000000000000001100110100001", -- 6560 FREE #<CONS 0 6561>
 "00000000000000000001100110100010", -- 6561 FREE #<CONS 0 6562>
 "00000000000000000001100110100011", -- 6562 FREE #<CONS 0 6563>
 "00000000000000000001100110100100", -- 6563 FREE #<CONS 0 6564>
 "00000000000000000001100110100101", -- 6564 FREE #<CONS 0 6565>
 "00000000000000000001100110100110", -- 6565 FREE #<CONS 0 6566>
 "00000000000000000001100110100111", -- 6566 FREE #<CONS 0 6567>
 "00000000000000000001100110101000", -- 6567 FREE #<CONS 0 6568>
 "00000000000000000001100110101001", -- 6568 FREE #<CONS 0 6569>
 "00000000000000000001100110101010", -- 6569 FREE #<CONS 0 6570>
 "00000000000000000001100110101011", -- 6570 FREE #<CONS 0 6571>
 "00000000000000000001100110101100", -- 6571 FREE #<CONS 0 6572>
 "00000000000000000001100110101101", -- 6572 FREE #<CONS 0 6573>
 "00000000000000000001100110101110", -- 6573 FREE #<CONS 0 6574>
 "00000000000000000001100110101111", -- 6574 FREE #<CONS 0 6575>
 "00000000000000000001100110110000", -- 6575 FREE #<CONS 0 6576>
 "00000000000000000001100110110001", -- 6576 FREE #<CONS 0 6577>
 "00000000000000000001100110110010", -- 6577 FREE #<CONS 0 6578>
 "00000000000000000001100110110011", -- 6578 FREE #<CONS 0 6579>
 "00000000000000000001100110110100", -- 6579 FREE #<CONS 0 6580>
 "00000000000000000001100110110101", -- 6580 FREE #<CONS 0 6581>
 "00000000000000000001100110110110", -- 6581 FREE #<CONS 0 6582>
 "00000000000000000001100110110111", -- 6582 FREE #<CONS 0 6583>
 "00000000000000000001100110111000", -- 6583 FREE #<CONS 0 6584>
 "00000000000000000001100110111001", -- 6584 FREE #<CONS 0 6585>
 "00000000000000000001100110111010", -- 6585 FREE #<CONS 0 6586>
 "00000000000000000001100110111011", -- 6586 FREE #<CONS 0 6587>
 "00000000000000000001100110111100", -- 6587 FREE #<CONS 0 6588>
 "00000000000000000001100110111101", -- 6588 FREE #<CONS 0 6589>
 "00000000000000000001100110111110", -- 6589 FREE #<CONS 0 6590>
 "00000000000000000001100110111111", -- 6590 FREE #<CONS 0 6591>
 "00000000000000000001100111000000", -- 6591 FREE #<CONS 0 6592>
 "00000000000000000001100111000001", -- 6592 FREE #<CONS 0 6593>
 "00000000000000000001100111000010", -- 6593 FREE #<CONS 0 6594>
 "00000000000000000001100111000011", -- 6594 FREE #<CONS 0 6595>
 "00000000000000000001100111000100", -- 6595 FREE #<CONS 0 6596>
 "00000000000000000001100111000101", -- 6596 FREE #<CONS 0 6597>
 "00000000000000000001100111000110", -- 6597 FREE #<CONS 0 6598>
 "00000000000000000001100111000111", -- 6598 FREE #<CONS 0 6599>
 "00000000000000000001100111001000", -- 6599 FREE #<CONS 0 6600>
 "00000000000000000001100111001001", -- 6600 FREE #<CONS 0 6601>
 "00000000000000000001100111001010", -- 6601 FREE #<CONS 0 6602>
 "00000000000000000001100111001011", -- 6602 FREE #<CONS 0 6603>
 "00000000000000000001100111001100", -- 6603 FREE #<CONS 0 6604>
 "00000000000000000001100111001101", -- 6604 FREE #<CONS 0 6605>
 "00000000000000000001100111001110", -- 6605 FREE #<CONS 0 6606>
 "00000000000000000001100111001111", -- 6606 FREE #<CONS 0 6607>
 "00000000000000000001100111010000", -- 6607 FREE #<CONS 0 6608>
 "00000000000000000001100111010001", -- 6608 FREE #<CONS 0 6609>
 "00000000000000000001100111010010", -- 6609 FREE #<CONS 0 6610>
 "00000000000000000001100111010011", -- 6610 FREE #<CONS 0 6611>
 "00000000000000000001100111010100", -- 6611 FREE #<CONS 0 6612>
 "00000000000000000001100111010101", -- 6612 FREE #<CONS 0 6613>
 "00000000000000000001100111010110", -- 6613 FREE #<CONS 0 6614>
 "00000000000000000001100111010111", -- 6614 FREE #<CONS 0 6615>
 "00000000000000000001100111011000", -- 6615 FREE #<CONS 0 6616>
 "00000000000000000001100111011001", -- 6616 FREE #<CONS 0 6617>
 "00000000000000000001100111011010", -- 6617 FREE #<CONS 0 6618>
 "00000000000000000001100111011011", -- 6618 FREE #<CONS 0 6619>
 "00000000000000000001100111011100", -- 6619 FREE #<CONS 0 6620>
 "00000000000000000001100111011101", -- 6620 FREE #<CONS 0 6621>
 "00000000000000000001100111011110", -- 6621 FREE #<CONS 0 6622>
 "00000000000000000001100111011111", -- 6622 FREE #<CONS 0 6623>
 "00000000000000000001100111100000", -- 6623 FREE #<CONS 0 6624>
 "00000000000000000001100111100001", -- 6624 FREE #<CONS 0 6625>
 "00000000000000000001100111100010", -- 6625 FREE #<CONS 0 6626>
 "00000000000000000001100111100011", -- 6626 FREE #<CONS 0 6627>
 "00000000000000000001100111100100", -- 6627 FREE #<CONS 0 6628>
 "00000000000000000001100111100101", -- 6628 FREE #<CONS 0 6629>
 "00000000000000000001100111100110", -- 6629 FREE #<CONS 0 6630>
 "00000000000000000001100111100111", -- 6630 FREE #<CONS 0 6631>
 "00000000000000000001100111101000", -- 6631 FREE #<CONS 0 6632>
 "00000000000000000001100111101001", -- 6632 FREE #<CONS 0 6633>
 "00000000000000000001100111101010", -- 6633 FREE #<CONS 0 6634>
 "00000000000000000001100111101011", -- 6634 FREE #<CONS 0 6635>
 "00000000000000000001100111101100", -- 6635 FREE #<CONS 0 6636>
 "00000000000000000001100111101101", -- 6636 FREE #<CONS 0 6637>
 "00000000000000000001100111101110", -- 6637 FREE #<CONS 0 6638>
 "00000000000000000001100111101111", -- 6638 FREE #<CONS 0 6639>
 "00000000000000000001100111110000", -- 6639 FREE #<CONS 0 6640>
 "00000000000000000001100111110001", -- 6640 FREE #<CONS 0 6641>
 "00000000000000000001100111110010", -- 6641 FREE #<CONS 0 6642>
 "00000000000000000001100111110011", -- 6642 FREE #<CONS 0 6643>
 "00000000000000000001100111110100", -- 6643 FREE #<CONS 0 6644>
 "00000000000000000001100111110101", -- 6644 FREE #<CONS 0 6645>
 "00000000000000000001100111110110", -- 6645 FREE #<CONS 0 6646>
 "00000000000000000001100111110111", -- 6646 FREE #<CONS 0 6647>
 "00000000000000000001100111111000", -- 6647 FREE #<CONS 0 6648>
 "00000000000000000001100111111001", -- 6648 FREE #<CONS 0 6649>
 "00000000000000000001100111111010", -- 6649 FREE #<CONS 0 6650>
 "00000000000000000001100111111011", -- 6650 FREE #<CONS 0 6651>
 "00000000000000000001100111111100", -- 6651 FREE #<CONS 0 6652>
 "00000000000000000001100111111101", -- 6652 FREE #<CONS 0 6653>
 "00000000000000000001100111111110", -- 6653 FREE #<CONS 0 6654>
 "00000000000000000001100111111111", -- 6654 FREE #<CONS 0 6655>
 "00000000000000000001101000000000", -- 6655 FREE #<CONS 0 6656>
 "00000000000000000001101000000001", -- 6656 FREE #<CONS 0 6657>
 "00000000000000000001101000000010", -- 6657 FREE #<CONS 0 6658>
 "00000000000000000001101000000011", -- 6658 FREE #<CONS 0 6659>
 "00000000000000000001101000000100", -- 6659 FREE #<CONS 0 6660>
 "00000000000000000001101000000101", -- 6660 FREE #<CONS 0 6661>
 "00000000000000000001101000000110", -- 6661 FREE #<CONS 0 6662>
 "00000000000000000001101000000111", -- 6662 FREE #<CONS 0 6663>
 "00000000000000000001101000001000", -- 6663 FREE #<CONS 0 6664>
 "00000000000000000001101000001001", -- 6664 FREE #<CONS 0 6665>
 "00000000000000000001101000001010", -- 6665 FREE #<CONS 0 6666>
 "00000000000000000001101000001011", -- 6666 FREE #<CONS 0 6667>
 "00000000000000000001101000001100", -- 6667 FREE #<CONS 0 6668>
 "00000000000000000001101000001101", -- 6668 FREE #<CONS 0 6669>
 "00000000000000000001101000001110", -- 6669 FREE #<CONS 0 6670>
 "00000000000000000001101000001111", -- 6670 FREE #<CONS 0 6671>
 "00000000000000000001101000010000", -- 6671 FREE #<CONS 0 6672>
 "00000000000000000001101000010001", -- 6672 FREE #<CONS 0 6673>
 "00000000000000000001101000010010", -- 6673 FREE #<CONS 0 6674>
 "00000000000000000001101000010011", -- 6674 FREE #<CONS 0 6675>
 "00000000000000000001101000010100", -- 6675 FREE #<CONS 0 6676>
 "00000000000000000001101000010101", -- 6676 FREE #<CONS 0 6677>
 "00000000000000000001101000010110", -- 6677 FREE #<CONS 0 6678>
 "00000000000000000001101000010111", -- 6678 FREE #<CONS 0 6679>
 "00000000000000000001101000011000", -- 6679 FREE #<CONS 0 6680>
 "00000000000000000001101000011001", -- 6680 FREE #<CONS 0 6681>
 "00000000000000000001101000011010", -- 6681 FREE #<CONS 0 6682>
 "00000000000000000001101000011011", -- 6682 FREE #<CONS 0 6683>
 "00000000000000000001101000011100", -- 6683 FREE #<CONS 0 6684>
 "00000000000000000001101000011101", -- 6684 FREE #<CONS 0 6685>
 "00000000000000000001101000011110", -- 6685 FREE #<CONS 0 6686>
 "00000000000000000001101000011111", -- 6686 FREE #<CONS 0 6687>
 "00000000000000000001101000100000", -- 6687 FREE #<CONS 0 6688>
 "00000000000000000001101000100001", -- 6688 FREE #<CONS 0 6689>
 "00000000000000000001101000100010", -- 6689 FREE #<CONS 0 6690>
 "00000000000000000001101000100011", -- 6690 FREE #<CONS 0 6691>
 "00000000000000000001101000100100", -- 6691 FREE #<CONS 0 6692>
 "00000000000000000001101000100101", -- 6692 FREE #<CONS 0 6693>
 "00000000000000000001101000100110", -- 6693 FREE #<CONS 0 6694>
 "00000000000000000001101000100111", -- 6694 FREE #<CONS 0 6695>
 "00000000000000000001101000101000", -- 6695 FREE #<CONS 0 6696>
 "00000000000000000001101000101001", -- 6696 FREE #<CONS 0 6697>
 "00000000000000000001101000101010", -- 6697 FREE #<CONS 0 6698>
 "00000000000000000001101000101011", -- 6698 FREE #<CONS 0 6699>
 "00000000000000000001101000101100", -- 6699 FREE #<CONS 0 6700>
 "00000000000000000001101000101101", -- 6700 FREE #<CONS 0 6701>
 "00000000000000000001101000101110", -- 6701 FREE #<CONS 0 6702>
 "00000000000000000001101000101111", -- 6702 FREE #<CONS 0 6703>
 "00000000000000000001101000110000", -- 6703 FREE #<CONS 0 6704>
 "00000000000000000001101000110001", -- 6704 FREE #<CONS 0 6705>
 "00000000000000000001101000110010", -- 6705 FREE #<CONS 0 6706>
 "00000000000000000001101000110011", -- 6706 FREE #<CONS 0 6707>
 "00000000000000000001101000110100", -- 6707 FREE #<CONS 0 6708>
 "00000000000000000001101000110101", -- 6708 FREE #<CONS 0 6709>
 "00000000000000000001101000110110", -- 6709 FREE #<CONS 0 6710>
 "00000000000000000001101000110111", -- 6710 FREE #<CONS 0 6711>
 "00000000000000000001101000111000", -- 6711 FREE #<CONS 0 6712>
 "00000000000000000001101000111001", -- 6712 FREE #<CONS 0 6713>
 "00000000000000000001101000111010", -- 6713 FREE #<CONS 0 6714>
 "00000000000000000001101000111011", -- 6714 FREE #<CONS 0 6715>
 "00000000000000000001101000111100", -- 6715 FREE #<CONS 0 6716>
 "00000000000000000001101000111101", -- 6716 FREE #<CONS 0 6717>
 "00000000000000000001101000111110", -- 6717 FREE #<CONS 0 6718>
 "00000000000000000001101000111111", -- 6718 FREE #<CONS 0 6719>
 "00000000000000000001101001000000", -- 6719 FREE #<CONS 0 6720>
 "00000000000000000001101001000001", -- 6720 FREE #<CONS 0 6721>
 "00000000000000000001101001000010", -- 6721 FREE #<CONS 0 6722>
 "00000000000000000001101001000011", -- 6722 FREE #<CONS 0 6723>
 "00000000000000000001101001000100", -- 6723 FREE #<CONS 0 6724>
 "00000000000000000001101001000101", -- 6724 FREE #<CONS 0 6725>
 "00000000000000000001101001000110", -- 6725 FREE #<CONS 0 6726>
 "00000000000000000001101001000111", -- 6726 FREE #<CONS 0 6727>
 "00000000000000000001101001001000", -- 6727 FREE #<CONS 0 6728>
 "00000000000000000001101001001001", -- 6728 FREE #<CONS 0 6729>
 "00000000000000000001101001001010", -- 6729 FREE #<CONS 0 6730>
 "00000000000000000001101001001011", -- 6730 FREE #<CONS 0 6731>
 "00000000000000000001101001001100", -- 6731 FREE #<CONS 0 6732>
 "00000000000000000001101001001101", -- 6732 FREE #<CONS 0 6733>
 "00000000000000000001101001001110", -- 6733 FREE #<CONS 0 6734>
 "00000000000000000001101001001111", -- 6734 FREE #<CONS 0 6735>
 "00000000000000000001101001010000", -- 6735 FREE #<CONS 0 6736>
 "00000000000000000001101001010001", -- 6736 FREE #<CONS 0 6737>
 "00000000000000000001101001010010", -- 6737 FREE #<CONS 0 6738>
 "00000000000000000001101001010011", -- 6738 FREE #<CONS 0 6739>
 "00000000000000000001101001010100", -- 6739 FREE #<CONS 0 6740>
 "00000000000000000001101001010101", -- 6740 FREE #<CONS 0 6741>
 "00000000000000000001101001010110", -- 6741 FREE #<CONS 0 6742>
 "00000000000000000001101001010111", -- 6742 FREE #<CONS 0 6743>
 "00000000000000000001101001011000", -- 6743 FREE #<CONS 0 6744>
 "00000000000000000001101001011001", -- 6744 FREE #<CONS 0 6745>
 "00000000000000000001101001011010", -- 6745 FREE #<CONS 0 6746>
 "00000000000000000001101001011011", -- 6746 FREE #<CONS 0 6747>
 "00000000000000000001101001011100", -- 6747 FREE #<CONS 0 6748>
 "00000000000000000001101001011101", -- 6748 FREE #<CONS 0 6749>
 "00000000000000000001101001011110", -- 6749 FREE #<CONS 0 6750>
 "00000000000000000001101001011111", -- 6750 FREE #<CONS 0 6751>
 "00000000000000000001101001100000", -- 6751 FREE #<CONS 0 6752>
 "00000000000000000001101001100001", -- 6752 FREE #<CONS 0 6753>
 "00000000000000000001101001100010", -- 6753 FREE #<CONS 0 6754>
 "00000000000000000001101001100011", -- 6754 FREE #<CONS 0 6755>
 "00000000000000000001101001100100", -- 6755 FREE #<CONS 0 6756>
 "00000000000000000001101001100101", -- 6756 FREE #<CONS 0 6757>
 "00000000000000000001101001100110", -- 6757 FREE #<CONS 0 6758>
 "00000000000000000001101001100111", -- 6758 FREE #<CONS 0 6759>
 "00000000000000000001101001101000", -- 6759 FREE #<CONS 0 6760>
 "00000000000000000001101001101001", -- 6760 FREE #<CONS 0 6761>
 "00000000000000000001101001101010", -- 6761 FREE #<CONS 0 6762>
 "00000000000000000001101001101011", -- 6762 FREE #<CONS 0 6763>
 "00000000000000000001101001101100", -- 6763 FREE #<CONS 0 6764>
 "00000000000000000001101001101101", -- 6764 FREE #<CONS 0 6765>
 "00000000000000000001101001101110", -- 6765 FREE #<CONS 0 6766>
 "00000000000000000001101001101111", -- 6766 FREE #<CONS 0 6767>
 "00000000000000000001101001110000", -- 6767 FREE #<CONS 0 6768>
 "00000000000000000001101001110001", -- 6768 FREE #<CONS 0 6769>
 "00000000000000000001101001110010", -- 6769 FREE #<CONS 0 6770>
 "00000000000000000001101001110011", -- 6770 FREE #<CONS 0 6771>
 "00000000000000000001101001110100", -- 6771 FREE #<CONS 0 6772>
 "00000000000000000001101001110101", -- 6772 FREE #<CONS 0 6773>
 "00000000000000000001101001110110", -- 6773 FREE #<CONS 0 6774>
 "00000000000000000001101001110111", -- 6774 FREE #<CONS 0 6775>
 "00000000000000000001101001111000", -- 6775 FREE #<CONS 0 6776>
 "00000000000000000001101001111001", -- 6776 FREE #<CONS 0 6777>
 "00000000000000000001101001111010", -- 6777 FREE #<CONS 0 6778>
 "00000000000000000001101001111011", -- 6778 FREE #<CONS 0 6779>
 "00000000000000000001101001111100", -- 6779 FREE #<CONS 0 6780>
 "00000000000000000001101001111101", -- 6780 FREE #<CONS 0 6781>
 "00000000000000000001101001111110", -- 6781 FREE #<CONS 0 6782>
 "00000000000000000001101001111111", -- 6782 FREE #<CONS 0 6783>
 "00000000000000000001101010000000", -- 6783 FREE #<CONS 0 6784>
 "00000000000000000001101010000001", -- 6784 FREE #<CONS 0 6785>
 "00000000000000000001101010000010", -- 6785 FREE #<CONS 0 6786>
 "00000000000000000001101010000011", -- 6786 FREE #<CONS 0 6787>
 "00000000000000000001101010000100", -- 6787 FREE #<CONS 0 6788>
 "00000000000000000001101010000101", -- 6788 FREE #<CONS 0 6789>
 "00000000000000000001101010000110", -- 6789 FREE #<CONS 0 6790>
 "00000000000000000001101010000111", -- 6790 FREE #<CONS 0 6791>
 "00000000000000000001101010001000", -- 6791 FREE #<CONS 0 6792>
 "00000000000000000001101010001001", -- 6792 FREE #<CONS 0 6793>
 "00000000000000000001101010001010", -- 6793 FREE #<CONS 0 6794>
 "00000000000000000001101010001011", -- 6794 FREE #<CONS 0 6795>
 "00000000000000000001101010001100", -- 6795 FREE #<CONS 0 6796>
 "00000000000000000001101010001101", -- 6796 FREE #<CONS 0 6797>
 "00000000000000000001101010001110", -- 6797 FREE #<CONS 0 6798>
 "00000000000000000001101010001111", -- 6798 FREE #<CONS 0 6799>
 "00000000000000000001101010010000", -- 6799 FREE #<CONS 0 6800>
 "00000000000000000001101010010001", -- 6800 FREE #<CONS 0 6801>
 "00000000000000000001101010010010", -- 6801 FREE #<CONS 0 6802>
 "00000000000000000001101010010011", -- 6802 FREE #<CONS 0 6803>
 "00000000000000000001101010010100", -- 6803 FREE #<CONS 0 6804>
 "00000000000000000001101010010101", -- 6804 FREE #<CONS 0 6805>
 "00000000000000000001101010010110", -- 6805 FREE #<CONS 0 6806>
 "00000000000000000001101010010111", -- 6806 FREE #<CONS 0 6807>
 "00000000000000000001101010011000", -- 6807 FREE #<CONS 0 6808>
 "00000000000000000001101010011001", -- 6808 FREE #<CONS 0 6809>
 "00000000000000000001101010011010", -- 6809 FREE #<CONS 0 6810>
 "00000000000000000001101010011011", -- 6810 FREE #<CONS 0 6811>
 "00000000000000000001101010011100", -- 6811 FREE #<CONS 0 6812>
 "00000000000000000001101010011101", -- 6812 FREE #<CONS 0 6813>
 "00000000000000000001101010011110", -- 6813 FREE #<CONS 0 6814>
 "00000000000000000001101010011111", -- 6814 FREE #<CONS 0 6815>
 "00000000000000000001101010100000", -- 6815 FREE #<CONS 0 6816>
 "00000000000000000001101010100001", -- 6816 FREE #<CONS 0 6817>
 "00000000000000000001101010100010", -- 6817 FREE #<CONS 0 6818>
 "00000000000000000001101010100011", -- 6818 FREE #<CONS 0 6819>
 "00000000000000000001101010100100", -- 6819 FREE #<CONS 0 6820>
 "00000000000000000001101010100101", -- 6820 FREE #<CONS 0 6821>
 "00000000000000000001101010100110", -- 6821 FREE #<CONS 0 6822>
 "00000000000000000001101010100111", -- 6822 FREE #<CONS 0 6823>
 "00000000000000000001101010101000", -- 6823 FREE #<CONS 0 6824>
 "00000000000000000001101010101001", -- 6824 FREE #<CONS 0 6825>
 "00000000000000000001101010101010", -- 6825 FREE #<CONS 0 6826>
 "00000000000000000001101010101011", -- 6826 FREE #<CONS 0 6827>
 "00000000000000000001101010101100", -- 6827 FREE #<CONS 0 6828>
 "00000000000000000001101010101101", -- 6828 FREE #<CONS 0 6829>
 "00000000000000000001101010101110", -- 6829 FREE #<CONS 0 6830>
 "00000000000000000001101010101111", -- 6830 FREE #<CONS 0 6831>
 "00000000000000000001101010110000", -- 6831 FREE #<CONS 0 6832>
 "00000000000000000001101010110001", -- 6832 FREE #<CONS 0 6833>
 "00000000000000000001101010110010", -- 6833 FREE #<CONS 0 6834>
 "00000000000000000001101010110011", -- 6834 FREE #<CONS 0 6835>
 "00000000000000000001101010110100", -- 6835 FREE #<CONS 0 6836>
 "00000000000000000001101010110101", -- 6836 FREE #<CONS 0 6837>
 "00000000000000000001101010110110", -- 6837 FREE #<CONS 0 6838>
 "00000000000000000001101010110111", -- 6838 FREE #<CONS 0 6839>
 "00000000000000000001101010111000", -- 6839 FREE #<CONS 0 6840>
 "00000000000000000001101010111001", -- 6840 FREE #<CONS 0 6841>
 "00000000000000000001101010111010", -- 6841 FREE #<CONS 0 6842>
 "00000000000000000001101010111011", -- 6842 FREE #<CONS 0 6843>
 "00000000000000000001101010111100", -- 6843 FREE #<CONS 0 6844>
 "00000000000000000001101010111101", -- 6844 FREE #<CONS 0 6845>
 "00000000000000000001101010111110", -- 6845 FREE #<CONS 0 6846>
 "00000000000000000001101010111111", -- 6846 FREE #<CONS 0 6847>
 "00000000000000000001101011000000", -- 6847 FREE #<CONS 0 6848>
 "00000000000000000001101011000001", -- 6848 FREE #<CONS 0 6849>
 "00000000000000000001101011000010", -- 6849 FREE #<CONS 0 6850>
 "00000000000000000001101011000011", -- 6850 FREE #<CONS 0 6851>
 "00000000000000000001101011000100", -- 6851 FREE #<CONS 0 6852>
 "00000000000000000001101011000101", -- 6852 FREE #<CONS 0 6853>
 "00000000000000000001101011000110", -- 6853 FREE #<CONS 0 6854>
 "00000000000000000001101011000111", -- 6854 FREE #<CONS 0 6855>
 "00000000000000000001101011001000", -- 6855 FREE #<CONS 0 6856>
 "00000000000000000001101011001001", -- 6856 FREE #<CONS 0 6857>
 "00000000000000000001101011001010", -- 6857 FREE #<CONS 0 6858>
 "00000000000000000001101011001011", -- 6858 FREE #<CONS 0 6859>
 "00000000000000000001101011001100", -- 6859 FREE #<CONS 0 6860>
 "00000000000000000001101011001101", -- 6860 FREE #<CONS 0 6861>
 "00000000000000000001101011001110", -- 6861 FREE #<CONS 0 6862>
 "00000000000000000001101011001111", -- 6862 FREE #<CONS 0 6863>
 "00000000000000000001101011010000", -- 6863 FREE #<CONS 0 6864>
 "00000000000000000001101011010001", -- 6864 FREE #<CONS 0 6865>
 "00000000000000000001101011010010", -- 6865 FREE #<CONS 0 6866>
 "00000000000000000001101011010011", -- 6866 FREE #<CONS 0 6867>
 "00000000000000000001101011010100", -- 6867 FREE #<CONS 0 6868>
 "00000000000000000001101011010101", -- 6868 FREE #<CONS 0 6869>
 "00000000000000000001101011010110", -- 6869 FREE #<CONS 0 6870>
 "00000000000000000001101011010111", -- 6870 FREE #<CONS 0 6871>
 "00000000000000000001101011011000", -- 6871 FREE #<CONS 0 6872>
 "00000000000000000001101011011001", -- 6872 FREE #<CONS 0 6873>
 "00000000000000000001101011011010", -- 6873 FREE #<CONS 0 6874>
 "00000000000000000001101011011011", -- 6874 FREE #<CONS 0 6875>
 "00000000000000000001101011011100", -- 6875 FREE #<CONS 0 6876>
 "00000000000000000001101011011101", -- 6876 FREE #<CONS 0 6877>
 "00000000000000000001101011011110", -- 6877 FREE #<CONS 0 6878>
 "00000000000000000001101011011111", -- 6878 FREE #<CONS 0 6879>
 "00000000000000000001101011100000", -- 6879 FREE #<CONS 0 6880>
 "00000000000000000001101011100001", -- 6880 FREE #<CONS 0 6881>
 "00000000000000000001101011100010", -- 6881 FREE #<CONS 0 6882>
 "00000000000000000001101011100011", -- 6882 FREE #<CONS 0 6883>
 "00000000000000000001101011100100", -- 6883 FREE #<CONS 0 6884>
 "00000000000000000001101011100101", -- 6884 FREE #<CONS 0 6885>
 "00000000000000000001101011100110", -- 6885 FREE #<CONS 0 6886>
 "00000000000000000001101011100111", -- 6886 FREE #<CONS 0 6887>
 "00000000000000000001101011101000", -- 6887 FREE #<CONS 0 6888>
 "00000000000000000001101011101001", -- 6888 FREE #<CONS 0 6889>
 "00000000000000000001101011101010", -- 6889 FREE #<CONS 0 6890>
 "00000000000000000001101011101011", -- 6890 FREE #<CONS 0 6891>
 "00000000000000000001101011101100", -- 6891 FREE #<CONS 0 6892>
 "00000000000000000001101011101101", -- 6892 FREE #<CONS 0 6893>
 "00000000000000000001101011101110", -- 6893 FREE #<CONS 0 6894>
 "00000000000000000001101011101111", -- 6894 FREE #<CONS 0 6895>
 "00000000000000000001101011110000", -- 6895 FREE #<CONS 0 6896>
 "00000000000000000001101011110001", -- 6896 FREE #<CONS 0 6897>
 "00000000000000000001101011110010", -- 6897 FREE #<CONS 0 6898>
 "00000000000000000001101011110011", -- 6898 FREE #<CONS 0 6899>
 "00000000000000000001101011110100", -- 6899 FREE #<CONS 0 6900>
 "00000000000000000001101011110101", -- 6900 FREE #<CONS 0 6901>
 "00000000000000000001101011110110", -- 6901 FREE #<CONS 0 6902>
 "00000000000000000001101011110111", -- 6902 FREE #<CONS 0 6903>
 "00000000000000000001101011111000", -- 6903 FREE #<CONS 0 6904>
 "00000000000000000001101011111001", -- 6904 FREE #<CONS 0 6905>
 "00000000000000000001101011111010", -- 6905 FREE #<CONS 0 6906>
 "00000000000000000001101011111011", -- 6906 FREE #<CONS 0 6907>
 "00000000000000000001101011111100", -- 6907 FREE #<CONS 0 6908>
 "00000000000000000001101011111101", -- 6908 FREE #<CONS 0 6909>
 "00000000000000000001101011111110", -- 6909 FREE #<CONS 0 6910>
 "00000000000000000001101011111111", -- 6910 FREE #<CONS 0 6911>
 "00000000000000000001101100000000", -- 6911 FREE #<CONS 0 6912>
 "00000000000000000001101100000001", -- 6912 FREE #<CONS 0 6913>
 "00000000000000000001101100000010", -- 6913 FREE #<CONS 0 6914>
 "00000000000000000001101100000011", -- 6914 FREE #<CONS 0 6915>
 "00000000000000000001101100000100", -- 6915 FREE #<CONS 0 6916>
 "00000000000000000001101100000101", -- 6916 FREE #<CONS 0 6917>
 "00000000000000000001101100000110", -- 6917 FREE #<CONS 0 6918>
 "00000000000000000001101100000111", -- 6918 FREE #<CONS 0 6919>
 "00000000000000000001101100001000", -- 6919 FREE #<CONS 0 6920>
 "00000000000000000001101100001001", -- 6920 FREE #<CONS 0 6921>
 "00000000000000000001101100001010", -- 6921 FREE #<CONS 0 6922>
 "00000000000000000001101100001011", -- 6922 FREE #<CONS 0 6923>
 "00000000000000000001101100001100", -- 6923 FREE #<CONS 0 6924>
 "00000000000000000001101100001101", -- 6924 FREE #<CONS 0 6925>
 "00000000000000000001101100001110", -- 6925 FREE #<CONS 0 6926>
 "00000000000000000001101100001111", -- 6926 FREE #<CONS 0 6927>
 "00000000000000000001101100010000", -- 6927 FREE #<CONS 0 6928>
 "00000000000000000001101100010001", -- 6928 FREE #<CONS 0 6929>
 "00000000000000000001101100010010", -- 6929 FREE #<CONS 0 6930>
 "00000000000000000001101100010011", -- 6930 FREE #<CONS 0 6931>
 "00000000000000000001101100010100", -- 6931 FREE #<CONS 0 6932>
 "00000000000000000001101100010101", -- 6932 FREE #<CONS 0 6933>
 "00000000000000000001101100010110", -- 6933 FREE #<CONS 0 6934>
 "00000000000000000001101100010111", -- 6934 FREE #<CONS 0 6935>
 "00000000000000000001101100011000", -- 6935 FREE #<CONS 0 6936>
 "00000000000000000001101100011001", -- 6936 FREE #<CONS 0 6937>
 "00000000000000000001101100011010", -- 6937 FREE #<CONS 0 6938>
 "00000000000000000001101100011011", -- 6938 FREE #<CONS 0 6939>
 "00000000000000000001101100011100", -- 6939 FREE #<CONS 0 6940>
 "00000000000000000001101100011101", -- 6940 FREE #<CONS 0 6941>
 "00000000000000000001101100011110", -- 6941 FREE #<CONS 0 6942>
 "00000000000000000001101100011111", -- 6942 FREE #<CONS 0 6943>
 "00000000000000000001101100100000", -- 6943 FREE #<CONS 0 6944>
 "00000000000000000001101100100001", -- 6944 FREE #<CONS 0 6945>
 "00000000000000000001101100100010", -- 6945 FREE #<CONS 0 6946>
 "00000000000000000001101100100011", -- 6946 FREE #<CONS 0 6947>
 "00000000000000000001101100100100", -- 6947 FREE #<CONS 0 6948>
 "00000000000000000001101100100101", -- 6948 FREE #<CONS 0 6949>
 "00000000000000000001101100100110", -- 6949 FREE #<CONS 0 6950>
 "00000000000000000001101100100111", -- 6950 FREE #<CONS 0 6951>
 "00000000000000000001101100101000", -- 6951 FREE #<CONS 0 6952>
 "00000000000000000001101100101001", -- 6952 FREE #<CONS 0 6953>
 "00000000000000000001101100101010", -- 6953 FREE #<CONS 0 6954>
 "00000000000000000001101100101011", -- 6954 FREE #<CONS 0 6955>
 "00000000000000000001101100101100", -- 6955 FREE #<CONS 0 6956>
 "00000000000000000001101100101101", -- 6956 FREE #<CONS 0 6957>
 "00000000000000000001101100101110", -- 6957 FREE #<CONS 0 6958>
 "00000000000000000001101100101111", -- 6958 FREE #<CONS 0 6959>
 "00000000000000000001101100110000", -- 6959 FREE #<CONS 0 6960>
 "00000000000000000001101100110001", -- 6960 FREE #<CONS 0 6961>
 "00000000000000000001101100110010", -- 6961 FREE #<CONS 0 6962>
 "00000000000000000001101100110011", -- 6962 FREE #<CONS 0 6963>
 "00000000000000000001101100110100", -- 6963 FREE #<CONS 0 6964>
 "00000000000000000001101100110101", -- 6964 FREE #<CONS 0 6965>
 "00000000000000000001101100110110", -- 6965 FREE #<CONS 0 6966>
 "00000000000000000001101100110111", -- 6966 FREE #<CONS 0 6967>
 "00000000000000000001101100111000", -- 6967 FREE #<CONS 0 6968>
 "00000000000000000001101100111001", -- 6968 FREE #<CONS 0 6969>
 "00000000000000000001101100111010", -- 6969 FREE #<CONS 0 6970>
 "00000000000000000001101100111011", -- 6970 FREE #<CONS 0 6971>
 "00000000000000000001101100111100", -- 6971 FREE #<CONS 0 6972>
 "00000000000000000001101100111101", -- 6972 FREE #<CONS 0 6973>
 "00000000000000000001101100111110", -- 6973 FREE #<CONS 0 6974>
 "00000000000000000001101100111111", -- 6974 FREE #<CONS 0 6975>
 "00000000000000000001101101000000", -- 6975 FREE #<CONS 0 6976>
 "00000000000000000001101101000001", -- 6976 FREE #<CONS 0 6977>
 "00000000000000000001101101000010", -- 6977 FREE #<CONS 0 6978>
 "00000000000000000001101101000011", -- 6978 FREE #<CONS 0 6979>
 "00000000000000000001101101000100", -- 6979 FREE #<CONS 0 6980>
 "00000000000000000001101101000101", -- 6980 FREE #<CONS 0 6981>
 "00000000000000000001101101000110", -- 6981 FREE #<CONS 0 6982>
 "00000000000000000001101101000111", -- 6982 FREE #<CONS 0 6983>
 "00000000000000000001101101001000", -- 6983 FREE #<CONS 0 6984>
 "00000000000000000001101101001001", -- 6984 FREE #<CONS 0 6985>
 "00000000000000000001101101001010", -- 6985 FREE #<CONS 0 6986>
 "00000000000000000001101101001011", -- 6986 FREE #<CONS 0 6987>
 "00000000000000000001101101001100", -- 6987 FREE #<CONS 0 6988>
 "00000000000000000001101101001101", -- 6988 FREE #<CONS 0 6989>
 "00000000000000000001101101001110", -- 6989 FREE #<CONS 0 6990>
 "00000000000000000001101101001111", -- 6990 FREE #<CONS 0 6991>
 "00000000000000000001101101010000", -- 6991 FREE #<CONS 0 6992>
 "00000000000000000001101101010001", -- 6992 FREE #<CONS 0 6993>
 "00000000000000000001101101010010", -- 6993 FREE #<CONS 0 6994>
 "00000000000000000001101101010011", -- 6994 FREE #<CONS 0 6995>
 "00000000000000000001101101010100", -- 6995 FREE #<CONS 0 6996>
 "00000000000000000001101101010101", -- 6996 FREE #<CONS 0 6997>
 "00000000000000000001101101010110", -- 6997 FREE #<CONS 0 6998>
 "00000000000000000001101101010111", -- 6998 FREE #<CONS 0 6999>
 "00000000000000000001101101011000", -- 6999 FREE #<CONS 0 7000>
 "00000000000000000001101101011001", -- 7000 FREE #<CONS 0 7001>
 "00000000000000000001101101011010", -- 7001 FREE #<CONS 0 7002>
 "00000000000000000001101101011011", -- 7002 FREE #<CONS 0 7003>
 "00000000000000000001101101011100", -- 7003 FREE #<CONS 0 7004>
 "00000000000000000001101101011101", -- 7004 FREE #<CONS 0 7005>
 "00000000000000000001101101011110", -- 7005 FREE #<CONS 0 7006>
 "00000000000000000001101101011111", -- 7006 FREE #<CONS 0 7007>
 "00000000000000000001101101100000", -- 7007 FREE #<CONS 0 7008>
 "00000000000000000001101101100001", -- 7008 FREE #<CONS 0 7009>
 "00000000000000000001101101100010", -- 7009 FREE #<CONS 0 7010>
 "00000000000000000001101101100011", -- 7010 FREE #<CONS 0 7011>
 "00000000000000000001101101100100", -- 7011 FREE #<CONS 0 7012>
 "00000000000000000001101101100101", -- 7012 FREE #<CONS 0 7013>
 "00000000000000000001101101100110", -- 7013 FREE #<CONS 0 7014>
 "00000000000000000001101101100111", -- 7014 FREE #<CONS 0 7015>
 "00000000000000000001101101101000", -- 7015 FREE #<CONS 0 7016>
 "00000000000000000001101101101001", -- 7016 FREE #<CONS 0 7017>
 "00000000000000000001101101101010", -- 7017 FREE #<CONS 0 7018>
 "00000000000000000001101101101011", -- 7018 FREE #<CONS 0 7019>
 "00000000000000000001101101101100", -- 7019 FREE #<CONS 0 7020>
 "00000000000000000001101101101101", -- 7020 FREE #<CONS 0 7021>
 "00000000000000000001101101101110", -- 7021 FREE #<CONS 0 7022>
 "00000000000000000001101101101111", -- 7022 FREE #<CONS 0 7023>
 "00000000000000000001101101110000", -- 7023 FREE #<CONS 0 7024>
 "00000000000000000001101101110001", -- 7024 FREE #<CONS 0 7025>
 "00000000000000000001101101110010", -- 7025 FREE #<CONS 0 7026>
 "00000000000000000001101101110011", -- 7026 FREE #<CONS 0 7027>
 "00000000000000000001101101110100", -- 7027 FREE #<CONS 0 7028>
 "00000000000000000001101101110101", -- 7028 FREE #<CONS 0 7029>
 "00000000000000000001101101110110", -- 7029 FREE #<CONS 0 7030>
 "00000000000000000001101101110111", -- 7030 FREE #<CONS 0 7031>
 "00000000000000000001101101111000", -- 7031 FREE #<CONS 0 7032>
 "00000000000000000001101101111001", -- 7032 FREE #<CONS 0 7033>
 "00000000000000000001101101111010", -- 7033 FREE #<CONS 0 7034>
 "00000000000000000001101101111011", -- 7034 FREE #<CONS 0 7035>
 "00000000000000000001101101111100", -- 7035 FREE #<CONS 0 7036>
 "00000000000000000001101101111101", -- 7036 FREE #<CONS 0 7037>
 "00000000000000000001101101111110", -- 7037 FREE #<CONS 0 7038>
 "00000000000000000001101101111111", -- 7038 FREE #<CONS 0 7039>
 "00000000000000000001101110000000", -- 7039 FREE #<CONS 0 7040>
 "00000000000000000001101110000001", -- 7040 FREE #<CONS 0 7041>
 "00000000000000000001101110000010", -- 7041 FREE #<CONS 0 7042>
 "00000000000000000001101110000011", -- 7042 FREE #<CONS 0 7043>
 "00000000000000000001101110000100", -- 7043 FREE #<CONS 0 7044>
 "00000000000000000001101110000101", -- 7044 FREE #<CONS 0 7045>
 "00000000000000000001101110000110", -- 7045 FREE #<CONS 0 7046>
 "00000000000000000001101110000111", -- 7046 FREE #<CONS 0 7047>
 "00000000000000000001101110001000", -- 7047 FREE #<CONS 0 7048>
 "00000000000000000001101110001001", -- 7048 FREE #<CONS 0 7049>
 "00000000000000000001101110001010", -- 7049 FREE #<CONS 0 7050>
 "00000000000000000001101110001011", -- 7050 FREE #<CONS 0 7051>
 "00000000000000000001101110001100", -- 7051 FREE #<CONS 0 7052>
 "00000000000000000001101110001101", -- 7052 FREE #<CONS 0 7053>
 "00000000000000000001101110001110", -- 7053 FREE #<CONS 0 7054>
 "00000000000000000001101110001111", -- 7054 FREE #<CONS 0 7055>
 "00000000000000000001101110010000", -- 7055 FREE #<CONS 0 7056>
 "00000000000000000001101110010001", -- 7056 FREE #<CONS 0 7057>
 "00000000000000000001101110010010", -- 7057 FREE #<CONS 0 7058>
 "00000000000000000001101110010011", -- 7058 FREE #<CONS 0 7059>
 "00000000000000000001101110010100", -- 7059 FREE #<CONS 0 7060>
 "00000000000000000001101110010101", -- 7060 FREE #<CONS 0 7061>
 "00000000000000000001101110010110", -- 7061 FREE #<CONS 0 7062>
 "00000000000000000001101110010111", -- 7062 FREE #<CONS 0 7063>
 "00000000000000000001101110011000", -- 7063 FREE #<CONS 0 7064>
 "00000000000000000001101110011001", -- 7064 FREE #<CONS 0 7065>
 "00000000000000000001101110011010", -- 7065 FREE #<CONS 0 7066>
 "00000000000000000001101110011011", -- 7066 FREE #<CONS 0 7067>
 "00000000000000000001101110011100", -- 7067 FREE #<CONS 0 7068>
 "00000000000000000001101110011101", -- 7068 FREE #<CONS 0 7069>
 "00000000000000000001101110011110", -- 7069 FREE #<CONS 0 7070>
 "00000000000000000001101110011111", -- 7070 FREE #<CONS 0 7071>
 "00000000000000000001101110100000", -- 7071 FREE #<CONS 0 7072>
 "00000000000000000001101110100001", -- 7072 FREE #<CONS 0 7073>
 "00000000000000000001101110100010", -- 7073 FREE #<CONS 0 7074>
 "00000000000000000001101110100011", -- 7074 FREE #<CONS 0 7075>
 "00000000000000000001101110100100", -- 7075 FREE #<CONS 0 7076>
 "00000000000000000001101110100101", -- 7076 FREE #<CONS 0 7077>
 "00000000000000000001101110100110", -- 7077 FREE #<CONS 0 7078>
 "00000000000000000001101110100111", -- 7078 FREE #<CONS 0 7079>
 "00000000000000000001101110101000", -- 7079 FREE #<CONS 0 7080>
 "00000000000000000001101110101001", -- 7080 FREE #<CONS 0 7081>
 "00000000000000000001101110101010", -- 7081 FREE #<CONS 0 7082>
 "00000000000000000001101110101011", -- 7082 FREE #<CONS 0 7083>
 "00000000000000000001101110101100", -- 7083 FREE #<CONS 0 7084>
 "00000000000000000001101110101101", -- 7084 FREE #<CONS 0 7085>
 "00000000000000000001101110101110", -- 7085 FREE #<CONS 0 7086>
 "00000000000000000001101110101111", -- 7086 FREE #<CONS 0 7087>
 "00000000000000000001101110110000", -- 7087 FREE #<CONS 0 7088>
 "00000000000000000001101110110001", -- 7088 FREE #<CONS 0 7089>
 "00000000000000000001101110110010", -- 7089 FREE #<CONS 0 7090>
 "00000000000000000001101110110011", -- 7090 FREE #<CONS 0 7091>
 "00000000000000000001101110110100", -- 7091 FREE #<CONS 0 7092>
 "00000000000000000001101110110101", -- 7092 FREE #<CONS 0 7093>
 "00000000000000000001101110110110", -- 7093 FREE #<CONS 0 7094>
 "00000000000000000001101110110111", -- 7094 FREE #<CONS 0 7095>
 "00000000000000000001101110111000", -- 7095 FREE #<CONS 0 7096>
 "00000000000000000001101110111001", -- 7096 FREE #<CONS 0 7097>
 "00000000000000000001101110111010", -- 7097 FREE #<CONS 0 7098>
 "00000000000000000001101110111011", -- 7098 FREE #<CONS 0 7099>
 "00000000000000000001101110111100", -- 7099 FREE #<CONS 0 7100>
 "00000000000000000001101110111101", -- 7100 FREE #<CONS 0 7101>
 "00000000000000000001101110111110", -- 7101 FREE #<CONS 0 7102>
 "00000000000000000001101110111111", -- 7102 FREE #<CONS 0 7103>
 "00000000000000000001101111000000", -- 7103 FREE #<CONS 0 7104>
 "00000000000000000001101111000001", -- 7104 FREE #<CONS 0 7105>
 "00000000000000000001101111000010", -- 7105 FREE #<CONS 0 7106>
 "00000000000000000001101111000011", -- 7106 FREE #<CONS 0 7107>
 "00000000000000000001101111000100", -- 7107 FREE #<CONS 0 7108>
 "00000000000000000001101111000101", -- 7108 FREE #<CONS 0 7109>
 "00000000000000000001101111000110", -- 7109 FREE #<CONS 0 7110>
 "00000000000000000001101111000111", -- 7110 FREE #<CONS 0 7111>
 "00000000000000000001101111001000", -- 7111 FREE #<CONS 0 7112>
 "00000000000000000001101111001001", -- 7112 FREE #<CONS 0 7113>
 "00000000000000000001101111001010", -- 7113 FREE #<CONS 0 7114>
 "00000000000000000001101111001011", -- 7114 FREE #<CONS 0 7115>
 "00000000000000000001101111001100", -- 7115 FREE #<CONS 0 7116>
 "00000000000000000001101111001101", -- 7116 FREE #<CONS 0 7117>
 "00000000000000000001101111001110", -- 7117 FREE #<CONS 0 7118>
 "00000000000000000001101111001111", -- 7118 FREE #<CONS 0 7119>
 "00000000000000000001101111010000", -- 7119 FREE #<CONS 0 7120>
 "00000000000000000001101111010001", -- 7120 FREE #<CONS 0 7121>
 "00000000000000000001101111010010", -- 7121 FREE #<CONS 0 7122>
 "00000000000000000001101111010011", -- 7122 FREE #<CONS 0 7123>
 "00000000000000000001101111010100", -- 7123 FREE #<CONS 0 7124>
 "00000000000000000001101111010101", -- 7124 FREE #<CONS 0 7125>
 "00000000000000000001101111010110", -- 7125 FREE #<CONS 0 7126>
 "00000000000000000001101111010111", -- 7126 FREE #<CONS 0 7127>
 "00000000000000000001101111011000", -- 7127 FREE #<CONS 0 7128>
 "00000000000000000001101111011001", -- 7128 FREE #<CONS 0 7129>
 "00000000000000000001101111011010", -- 7129 FREE #<CONS 0 7130>
 "00000000000000000001101111011011", -- 7130 FREE #<CONS 0 7131>
 "00000000000000000001101111011100", -- 7131 FREE #<CONS 0 7132>
 "00000000000000000001101111011101", -- 7132 FREE #<CONS 0 7133>
 "00000000000000000001101111011110", -- 7133 FREE #<CONS 0 7134>
 "00000000000000000001101111011111", -- 7134 FREE #<CONS 0 7135>
 "00000000000000000001101111100000", -- 7135 FREE #<CONS 0 7136>
 "00000000000000000001101111100001", -- 7136 FREE #<CONS 0 7137>
 "00000000000000000001101111100010", -- 7137 FREE #<CONS 0 7138>
 "00000000000000000001101111100011", -- 7138 FREE #<CONS 0 7139>
 "00000000000000000001101111100100", -- 7139 FREE #<CONS 0 7140>
 "00000000000000000001101111100101", -- 7140 FREE #<CONS 0 7141>
 "00000000000000000001101111100110", -- 7141 FREE #<CONS 0 7142>
 "00000000000000000001101111100111", -- 7142 FREE #<CONS 0 7143>
 "00000000000000000001101111101000", -- 7143 FREE #<CONS 0 7144>
 "00000000000000000001101111101001", -- 7144 FREE #<CONS 0 7145>
 "00000000000000000001101111101010", -- 7145 FREE #<CONS 0 7146>
 "00000000000000000001101111101011", -- 7146 FREE #<CONS 0 7147>
 "00000000000000000001101111101100", -- 7147 FREE #<CONS 0 7148>
 "00000000000000000001101111101101", -- 7148 FREE #<CONS 0 7149>
 "00000000000000000001101111101110", -- 7149 FREE #<CONS 0 7150>
 "00000000000000000001101111101111", -- 7150 FREE #<CONS 0 7151>
 "00000000000000000001101111110000", -- 7151 FREE #<CONS 0 7152>
 "00000000000000000001101111110001", -- 7152 FREE #<CONS 0 7153>
 "00000000000000000001101111110010", -- 7153 FREE #<CONS 0 7154>
 "00000000000000000001101111110011", -- 7154 FREE #<CONS 0 7155>
 "00000000000000000001101111110100", -- 7155 FREE #<CONS 0 7156>
 "00000000000000000001101111110101", -- 7156 FREE #<CONS 0 7157>
 "00000000000000000001101111110110", -- 7157 FREE #<CONS 0 7158>
 "00000000000000000001101111110111", -- 7158 FREE #<CONS 0 7159>
 "00000000000000000001101111111000", -- 7159 FREE #<CONS 0 7160>
 "00000000000000000001101111111001", -- 7160 FREE #<CONS 0 7161>
 "00000000000000000001101111111010", -- 7161 FREE #<CONS 0 7162>
 "00000000000000000001101111111011", -- 7162 FREE #<CONS 0 7163>
 "00000000000000000001101111111100", -- 7163 FREE #<CONS 0 7164>
 "00000000000000000001101111111101", -- 7164 FREE #<CONS 0 7165>
 "00000000000000000001101111111110", -- 7165 FREE #<CONS 0 7166>
 "00000000000000000001101111111111", -- 7166 FREE #<CONS 0 7167>
 "00000000000000000001110000000000", -- 7167 FREE #<CONS 0 7168>
 "00000000000000000001110000000001", -- 7168 FREE #<CONS 0 7169>
 "00000000000000000001110000000010", -- 7169 FREE #<CONS 0 7170>
 "00000000000000000001110000000011", -- 7170 FREE #<CONS 0 7171>
 "00000000000000000001110000000100", -- 7171 FREE #<CONS 0 7172>
 "00000000000000000001110000000101", -- 7172 FREE #<CONS 0 7173>
 "00000000000000000001110000000110", -- 7173 FREE #<CONS 0 7174>
 "00000000000000000001110000000111", -- 7174 FREE #<CONS 0 7175>
 "00000000000000000001110000001000", -- 7175 FREE #<CONS 0 7176>
 "00000000000000000001110000001001", -- 7176 FREE #<CONS 0 7177>
 "00000000000000000001110000001010", -- 7177 FREE #<CONS 0 7178>
 "00000000000000000001110000001011", -- 7178 FREE #<CONS 0 7179>
 "00000000000000000001110000001100", -- 7179 FREE #<CONS 0 7180>
 "00000000000000000001110000001101", -- 7180 FREE #<CONS 0 7181>
 "00000000000000000001110000001110", -- 7181 FREE #<CONS 0 7182>
 "00000000000000000001110000001111", -- 7182 FREE #<CONS 0 7183>
 "00000000000000000001110000010000", -- 7183 FREE #<CONS 0 7184>
 "00000000000000000001110000010001", -- 7184 FREE #<CONS 0 7185>
 "00000000000000000001110000010010", -- 7185 FREE #<CONS 0 7186>
 "00000000000000000001110000010011", -- 7186 FREE #<CONS 0 7187>
 "00000000000000000001110000010100", -- 7187 FREE #<CONS 0 7188>
 "00000000000000000001110000010101", -- 7188 FREE #<CONS 0 7189>
 "00000000000000000001110000010110", -- 7189 FREE #<CONS 0 7190>
 "00000000000000000001110000010111", -- 7190 FREE #<CONS 0 7191>
 "00000000000000000001110000011000", -- 7191 FREE #<CONS 0 7192>
 "00000000000000000001110000011001", -- 7192 FREE #<CONS 0 7193>
 "00000000000000000001110000011010", -- 7193 FREE #<CONS 0 7194>
 "00000000000000000001110000011011", -- 7194 FREE #<CONS 0 7195>
 "00000000000000000001110000011100", -- 7195 FREE #<CONS 0 7196>
 "00000000000000000001110000011101", -- 7196 FREE #<CONS 0 7197>
 "00000000000000000001110000011110", -- 7197 FREE #<CONS 0 7198>
 "00000000000000000001110000011111", -- 7198 FREE #<CONS 0 7199>
 "00000000000000000001110000100000", -- 7199 FREE #<CONS 0 7200>
 "00000000000000000001110000100001", -- 7200 FREE #<CONS 0 7201>
 "00000000000000000001110000100010", -- 7201 FREE #<CONS 0 7202>
 "00000000000000000001110000100011", -- 7202 FREE #<CONS 0 7203>
 "00000000000000000001110000100100", -- 7203 FREE #<CONS 0 7204>
 "00000000000000000001110000100101", -- 7204 FREE #<CONS 0 7205>
 "00000000000000000001110000100110", -- 7205 FREE #<CONS 0 7206>
 "00000000000000000001110000100111", -- 7206 FREE #<CONS 0 7207>
 "00000000000000000001110000101000", -- 7207 FREE #<CONS 0 7208>
 "00000000000000000001110000101001", -- 7208 FREE #<CONS 0 7209>
 "00000000000000000001110000101010", -- 7209 FREE #<CONS 0 7210>
 "00000000000000000001110000101011", -- 7210 FREE #<CONS 0 7211>
 "00000000000000000001110000101100", -- 7211 FREE #<CONS 0 7212>
 "00000000000000000001110000101101", -- 7212 FREE #<CONS 0 7213>
 "00000000000000000001110000101110", -- 7213 FREE #<CONS 0 7214>
 "00000000000000000001110000101111", -- 7214 FREE #<CONS 0 7215>
 "00000000000000000001110000110000", -- 7215 FREE #<CONS 0 7216>
 "00000000000000000001110000110001", -- 7216 FREE #<CONS 0 7217>
 "00000000000000000001110000110010", -- 7217 FREE #<CONS 0 7218>
 "00000000000000000001110000110011", -- 7218 FREE #<CONS 0 7219>
 "00000000000000000001110000110100", -- 7219 FREE #<CONS 0 7220>
 "00000000000000000001110000110101", -- 7220 FREE #<CONS 0 7221>
 "00000000000000000001110000110110", -- 7221 FREE #<CONS 0 7222>
 "00000000000000000001110000110111", -- 7222 FREE #<CONS 0 7223>
 "00000000000000000001110000111000", -- 7223 FREE #<CONS 0 7224>
 "00000000000000000001110000111001", -- 7224 FREE #<CONS 0 7225>
 "00000000000000000001110000111010", -- 7225 FREE #<CONS 0 7226>
 "00000000000000000001110000111011", -- 7226 FREE #<CONS 0 7227>
 "00000000000000000001110000111100", -- 7227 FREE #<CONS 0 7228>
 "00000000000000000001110000111101", -- 7228 FREE #<CONS 0 7229>
 "00000000000000000001110000111110", -- 7229 FREE #<CONS 0 7230>
 "00000000000000000001110000111111", -- 7230 FREE #<CONS 0 7231>
 "00000000000000000001110001000000", -- 7231 FREE #<CONS 0 7232>
 "00000000000000000001110001000001", -- 7232 FREE #<CONS 0 7233>
 "00000000000000000001110001000010", -- 7233 FREE #<CONS 0 7234>
 "00000000000000000001110001000011", -- 7234 FREE #<CONS 0 7235>
 "00000000000000000001110001000100", -- 7235 FREE #<CONS 0 7236>
 "00000000000000000001110001000101", -- 7236 FREE #<CONS 0 7237>
 "00000000000000000001110001000110", -- 7237 FREE #<CONS 0 7238>
 "00000000000000000001110001000111", -- 7238 FREE #<CONS 0 7239>
 "00000000000000000001110001001000", -- 7239 FREE #<CONS 0 7240>
 "00000000000000000001110001001001", -- 7240 FREE #<CONS 0 7241>
 "00000000000000000001110001001010", -- 7241 FREE #<CONS 0 7242>
 "00000000000000000001110001001011", -- 7242 FREE #<CONS 0 7243>
 "00000000000000000001110001001100", -- 7243 FREE #<CONS 0 7244>
 "00000000000000000001110001001101", -- 7244 FREE #<CONS 0 7245>
 "00000000000000000001110001001110", -- 7245 FREE #<CONS 0 7246>
 "00000000000000000001110001001111", -- 7246 FREE #<CONS 0 7247>
 "00000000000000000001110001010000", -- 7247 FREE #<CONS 0 7248>
 "00000000000000000001110001010001", -- 7248 FREE #<CONS 0 7249>
 "00000000000000000001110001010010", -- 7249 FREE #<CONS 0 7250>
 "00000000000000000001110001010011", -- 7250 FREE #<CONS 0 7251>
 "00000000000000000001110001010100", -- 7251 FREE #<CONS 0 7252>
 "00000000000000000001110001010101", -- 7252 FREE #<CONS 0 7253>
 "00000000000000000001110001010110", -- 7253 FREE #<CONS 0 7254>
 "00000000000000000001110001010111", -- 7254 FREE #<CONS 0 7255>
 "00000000000000000001110001011000", -- 7255 FREE #<CONS 0 7256>
 "00000000000000000001110001011001", -- 7256 FREE #<CONS 0 7257>
 "00000000000000000001110001011010", -- 7257 FREE #<CONS 0 7258>
 "00000000000000000001110001011011", -- 7258 FREE #<CONS 0 7259>
 "00000000000000000001110001011100", -- 7259 FREE #<CONS 0 7260>
 "00000000000000000001110001011101", -- 7260 FREE #<CONS 0 7261>
 "00000000000000000001110001011110", -- 7261 FREE #<CONS 0 7262>
 "00000000000000000001110001011111", -- 7262 FREE #<CONS 0 7263>
 "00000000000000000001110001100000", -- 7263 FREE #<CONS 0 7264>
 "00000000000000000001110001100001", -- 7264 FREE #<CONS 0 7265>
 "00000000000000000001110001100010", -- 7265 FREE #<CONS 0 7266>
 "00000000000000000001110001100011", -- 7266 FREE #<CONS 0 7267>
 "00000000000000000001110001100100", -- 7267 FREE #<CONS 0 7268>
 "00000000000000000001110001100101", -- 7268 FREE #<CONS 0 7269>
 "00000000000000000001110001100110", -- 7269 FREE #<CONS 0 7270>
 "00000000000000000001110001100111", -- 7270 FREE #<CONS 0 7271>
 "00000000000000000001110001101000", -- 7271 FREE #<CONS 0 7272>
 "00000000000000000001110001101001", -- 7272 FREE #<CONS 0 7273>
 "00000000000000000001110001101010", -- 7273 FREE #<CONS 0 7274>
 "00000000000000000001110001101011", -- 7274 FREE #<CONS 0 7275>
 "00000000000000000001110001101100", -- 7275 FREE #<CONS 0 7276>
 "00000000000000000001110001101101", -- 7276 FREE #<CONS 0 7277>
 "00000000000000000001110001101110", -- 7277 FREE #<CONS 0 7278>
 "00000000000000000001110001101111", -- 7278 FREE #<CONS 0 7279>
 "00000000000000000001110001110000", -- 7279 FREE #<CONS 0 7280>
 "00000000000000000001110001110001", -- 7280 FREE #<CONS 0 7281>
 "00000000000000000001110001110010", -- 7281 FREE #<CONS 0 7282>
 "00000000000000000001110001110011", -- 7282 FREE #<CONS 0 7283>
 "00000000000000000001110001110100", -- 7283 FREE #<CONS 0 7284>
 "00000000000000000001110001110101", -- 7284 FREE #<CONS 0 7285>
 "00000000000000000001110001110110", -- 7285 FREE #<CONS 0 7286>
 "00000000000000000001110001110111", -- 7286 FREE #<CONS 0 7287>
 "00000000000000000001110001111000", -- 7287 FREE #<CONS 0 7288>
 "00000000000000000001110001111001", -- 7288 FREE #<CONS 0 7289>
 "00000000000000000001110001111010", -- 7289 FREE #<CONS 0 7290>
 "00000000000000000001110001111011", -- 7290 FREE #<CONS 0 7291>
 "00000000000000000001110001111100", -- 7291 FREE #<CONS 0 7292>
 "00000000000000000001110001111101", -- 7292 FREE #<CONS 0 7293>
 "00000000000000000001110001111110", -- 7293 FREE #<CONS 0 7294>
 "00000000000000000001110001111111", -- 7294 FREE #<CONS 0 7295>
 "00000000000000000001110010000000", -- 7295 FREE #<CONS 0 7296>
 "00000000000000000001110010000001", -- 7296 FREE #<CONS 0 7297>
 "00000000000000000001110010000010", -- 7297 FREE #<CONS 0 7298>
 "00000000000000000001110010000011", -- 7298 FREE #<CONS 0 7299>
 "00000000000000000001110010000100", -- 7299 FREE #<CONS 0 7300>
 "00000000000000000001110010000101", -- 7300 FREE #<CONS 0 7301>
 "00000000000000000001110010000110", -- 7301 FREE #<CONS 0 7302>
 "00000000000000000001110010000111", -- 7302 FREE #<CONS 0 7303>
 "00000000000000000001110010001000", -- 7303 FREE #<CONS 0 7304>
 "00000000000000000001110010001001", -- 7304 FREE #<CONS 0 7305>
 "00000000000000000001110010001010", -- 7305 FREE #<CONS 0 7306>
 "00000000000000000001110010001011", -- 7306 FREE #<CONS 0 7307>
 "00000000000000000001110010001100", -- 7307 FREE #<CONS 0 7308>
 "00000000000000000001110010001101", -- 7308 FREE #<CONS 0 7309>
 "00000000000000000001110010001110", -- 7309 FREE #<CONS 0 7310>
 "00000000000000000001110010001111", -- 7310 FREE #<CONS 0 7311>
 "00000000000000000001110010010000", -- 7311 FREE #<CONS 0 7312>
 "00000000000000000001110010010001", -- 7312 FREE #<CONS 0 7313>
 "00000000000000000001110010010010", -- 7313 FREE #<CONS 0 7314>
 "00000000000000000001110010010011", -- 7314 FREE #<CONS 0 7315>
 "00000000000000000001110010010100", -- 7315 FREE #<CONS 0 7316>
 "00000000000000000001110010010101", -- 7316 FREE #<CONS 0 7317>
 "00000000000000000001110010010110", -- 7317 FREE #<CONS 0 7318>
 "00000000000000000001110010010111", -- 7318 FREE #<CONS 0 7319>
 "00000000000000000001110010011000", -- 7319 FREE #<CONS 0 7320>
 "00000000000000000001110010011001", -- 7320 FREE #<CONS 0 7321>
 "00000000000000000001110010011010", -- 7321 FREE #<CONS 0 7322>
 "00000000000000000001110010011011", -- 7322 FREE #<CONS 0 7323>
 "00000000000000000001110010011100", -- 7323 FREE #<CONS 0 7324>
 "00000000000000000001110010011101", -- 7324 FREE #<CONS 0 7325>
 "00000000000000000001110010011110", -- 7325 FREE #<CONS 0 7326>
 "00000000000000000001110010011111", -- 7326 FREE #<CONS 0 7327>
 "00000000000000000001110010100000", -- 7327 FREE #<CONS 0 7328>
 "00000000000000000001110010100001", -- 7328 FREE #<CONS 0 7329>
 "00000000000000000001110010100010", -- 7329 FREE #<CONS 0 7330>
 "00000000000000000001110010100011", -- 7330 FREE #<CONS 0 7331>
 "00000000000000000001110010100100", -- 7331 FREE #<CONS 0 7332>
 "00000000000000000001110010100101", -- 7332 FREE #<CONS 0 7333>
 "00000000000000000001110010100110", -- 7333 FREE #<CONS 0 7334>
 "00000000000000000001110010100111", -- 7334 FREE #<CONS 0 7335>
 "00000000000000000001110010101000", -- 7335 FREE #<CONS 0 7336>
 "00000000000000000001110010101001", -- 7336 FREE #<CONS 0 7337>
 "00000000000000000001110010101010", -- 7337 FREE #<CONS 0 7338>
 "00000000000000000001110010101011", -- 7338 FREE #<CONS 0 7339>
 "00000000000000000001110010101100", -- 7339 FREE #<CONS 0 7340>
 "00000000000000000001110010101101", -- 7340 FREE #<CONS 0 7341>
 "00000000000000000001110010101110", -- 7341 FREE #<CONS 0 7342>
 "00000000000000000001110010101111", -- 7342 FREE #<CONS 0 7343>
 "00000000000000000001110010110000", -- 7343 FREE #<CONS 0 7344>
 "00000000000000000001110010110001", -- 7344 FREE #<CONS 0 7345>
 "00000000000000000001110010110010", -- 7345 FREE #<CONS 0 7346>
 "00000000000000000001110010110011", -- 7346 FREE #<CONS 0 7347>
 "00000000000000000001110010110100", -- 7347 FREE #<CONS 0 7348>
 "00000000000000000001110010110101", -- 7348 FREE #<CONS 0 7349>
 "00000000000000000001110010110110", -- 7349 FREE #<CONS 0 7350>
 "00000000000000000001110010110111", -- 7350 FREE #<CONS 0 7351>
 "00000000000000000001110010111000", -- 7351 FREE #<CONS 0 7352>
 "00000000000000000001110010111001", -- 7352 FREE #<CONS 0 7353>
 "00000000000000000001110010111010", -- 7353 FREE #<CONS 0 7354>
 "00000000000000000001110010111011", -- 7354 FREE #<CONS 0 7355>
 "00000000000000000001110010111100", -- 7355 FREE #<CONS 0 7356>
 "00000000000000000001110010111101", -- 7356 FREE #<CONS 0 7357>
 "00000000000000000001110010111110", -- 7357 FREE #<CONS 0 7358>
 "00000000000000000001110010111111", -- 7358 FREE #<CONS 0 7359>
 "00000000000000000001110011000000", -- 7359 FREE #<CONS 0 7360>
 "00000000000000000001110011000001", -- 7360 FREE #<CONS 0 7361>
 "00000000000000000001110011000010", -- 7361 FREE #<CONS 0 7362>
 "00000000000000000001110011000011", -- 7362 FREE #<CONS 0 7363>
 "00000000000000000001110011000100", -- 7363 FREE #<CONS 0 7364>
 "00000000000000000001110011000101", -- 7364 FREE #<CONS 0 7365>
 "00000000000000000001110011000110", -- 7365 FREE #<CONS 0 7366>
 "00000000000000000001110011000111", -- 7366 FREE #<CONS 0 7367>
 "00000000000000000001110011001000", -- 7367 FREE #<CONS 0 7368>
 "00000000000000000001110011001001", -- 7368 FREE #<CONS 0 7369>
 "00000000000000000001110011001010", -- 7369 FREE #<CONS 0 7370>
 "00000000000000000001110011001011", -- 7370 FREE #<CONS 0 7371>
 "00000000000000000001110011001100", -- 7371 FREE #<CONS 0 7372>
 "00000000000000000001110011001101", -- 7372 FREE #<CONS 0 7373>
 "00000000000000000001110011001110", -- 7373 FREE #<CONS 0 7374>
 "00000000000000000001110011001111", -- 7374 FREE #<CONS 0 7375>
 "00000000000000000001110011010000", -- 7375 FREE #<CONS 0 7376>
 "00000000000000000001110011010001", -- 7376 FREE #<CONS 0 7377>
 "00000000000000000001110011010010", -- 7377 FREE #<CONS 0 7378>
 "00000000000000000001110011010011", -- 7378 FREE #<CONS 0 7379>
 "00000000000000000001110011010100", -- 7379 FREE #<CONS 0 7380>
 "00000000000000000001110011010101", -- 7380 FREE #<CONS 0 7381>
 "00000000000000000001110011010110", -- 7381 FREE #<CONS 0 7382>
 "00000000000000000001110011010111", -- 7382 FREE #<CONS 0 7383>
 "00000000000000000001110011011000", -- 7383 FREE #<CONS 0 7384>
 "00000000000000000001110011011001", -- 7384 FREE #<CONS 0 7385>
 "00000000000000000001110011011010", -- 7385 FREE #<CONS 0 7386>
 "00000000000000000001110011011011", -- 7386 FREE #<CONS 0 7387>
 "00000000000000000001110011011100", -- 7387 FREE #<CONS 0 7388>
 "00000000000000000001110011011101", -- 7388 FREE #<CONS 0 7389>
 "00000000000000000001110011011110", -- 7389 FREE #<CONS 0 7390>
 "00000000000000000001110011011111", -- 7390 FREE #<CONS 0 7391>
 "00000000000000000001110011100000", -- 7391 FREE #<CONS 0 7392>
 "00000000000000000001110011100001", -- 7392 FREE #<CONS 0 7393>
 "00000000000000000001110011100010", -- 7393 FREE #<CONS 0 7394>
 "00000000000000000001110011100011", -- 7394 FREE #<CONS 0 7395>
 "00000000000000000001110011100100", -- 7395 FREE #<CONS 0 7396>
 "00000000000000000001110011100101", -- 7396 FREE #<CONS 0 7397>
 "00000000000000000001110011100110", -- 7397 FREE #<CONS 0 7398>
 "00000000000000000001110011100111", -- 7398 FREE #<CONS 0 7399>
 "00000000000000000001110011101000", -- 7399 FREE #<CONS 0 7400>
 "00000000000000000001110011101001", -- 7400 FREE #<CONS 0 7401>
 "00000000000000000001110011101010", -- 7401 FREE #<CONS 0 7402>
 "00000000000000000001110011101011", -- 7402 FREE #<CONS 0 7403>
 "00000000000000000001110011101100", -- 7403 FREE #<CONS 0 7404>
 "00000000000000000001110011101101", -- 7404 FREE #<CONS 0 7405>
 "00000000000000000001110011101110", -- 7405 FREE #<CONS 0 7406>
 "00000000000000000001110011101111", -- 7406 FREE #<CONS 0 7407>
 "00000000000000000001110011110000", -- 7407 FREE #<CONS 0 7408>
 "00000000000000000001110011110001", -- 7408 FREE #<CONS 0 7409>
 "00000000000000000001110011110010", -- 7409 FREE #<CONS 0 7410>
 "00000000000000000001110011110011", -- 7410 FREE #<CONS 0 7411>
 "00000000000000000001110011110100", -- 7411 FREE #<CONS 0 7412>
 "00000000000000000001110011110101", -- 7412 FREE #<CONS 0 7413>
 "00000000000000000001110011110110", -- 7413 FREE #<CONS 0 7414>
 "00000000000000000001110011110111", -- 7414 FREE #<CONS 0 7415>
 "00000000000000000001110011111000", -- 7415 FREE #<CONS 0 7416>
 "00000000000000000001110011111001", -- 7416 FREE #<CONS 0 7417>
 "00000000000000000001110011111010", -- 7417 FREE #<CONS 0 7418>
 "00000000000000000001110011111011", -- 7418 FREE #<CONS 0 7419>
 "00000000000000000001110011111100", -- 7419 FREE #<CONS 0 7420>
 "00000000000000000001110011111101", -- 7420 FREE #<CONS 0 7421>
 "00000000000000000001110011111110", -- 7421 FREE #<CONS 0 7422>
 "00000000000000000001110011111111", -- 7422 FREE #<CONS 0 7423>
 "00000000000000000001110100000000", -- 7423 FREE #<CONS 0 7424>
 "00000000000000000001110100000001", -- 7424 FREE #<CONS 0 7425>
 "00000000000000000001110100000010", -- 7425 FREE #<CONS 0 7426>
 "00000000000000000001110100000011", -- 7426 FREE #<CONS 0 7427>
 "00000000000000000001110100000100", -- 7427 FREE #<CONS 0 7428>
 "00000000000000000001110100000101", -- 7428 FREE #<CONS 0 7429>
 "00000000000000000001110100000110", -- 7429 FREE #<CONS 0 7430>
 "00000000000000000001110100000111", -- 7430 FREE #<CONS 0 7431>
 "00000000000000000001110100001000", -- 7431 FREE #<CONS 0 7432>
 "00000000000000000001110100001001", -- 7432 FREE #<CONS 0 7433>
 "00000000000000000001110100001010", -- 7433 FREE #<CONS 0 7434>
 "00000000000000000001110100001011", -- 7434 FREE #<CONS 0 7435>
 "00000000000000000001110100001100", -- 7435 FREE #<CONS 0 7436>
 "00000000000000000001110100001101", -- 7436 FREE #<CONS 0 7437>
 "00000000000000000001110100001110", -- 7437 FREE #<CONS 0 7438>
 "00000000000000000001110100001111", -- 7438 FREE #<CONS 0 7439>
 "00000000000000000001110100010000", -- 7439 FREE #<CONS 0 7440>
 "00000000000000000001110100010001", -- 7440 FREE #<CONS 0 7441>
 "00000000000000000001110100010010", -- 7441 FREE #<CONS 0 7442>
 "00000000000000000001110100010011", -- 7442 FREE #<CONS 0 7443>
 "00000000000000000001110100010100", -- 7443 FREE #<CONS 0 7444>
 "00000000000000000001110100010101", -- 7444 FREE #<CONS 0 7445>
 "00000000000000000001110100010110", -- 7445 FREE #<CONS 0 7446>
 "00000000000000000001110100010111", -- 7446 FREE #<CONS 0 7447>
 "00000000000000000001110100011000", -- 7447 FREE #<CONS 0 7448>
 "00000000000000000001110100011001", -- 7448 FREE #<CONS 0 7449>
 "00000000000000000001110100011010", -- 7449 FREE #<CONS 0 7450>
 "00000000000000000001110100011011", -- 7450 FREE #<CONS 0 7451>
 "00000000000000000001110100011100", -- 7451 FREE #<CONS 0 7452>
 "00000000000000000001110100011101", -- 7452 FREE #<CONS 0 7453>
 "00000000000000000001110100011110", -- 7453 FREE #<CONS 0 7454>
 "00000000000000000001110100011111", -- 7454 FREE #<CONS 0 7455>
 "00000000000000000001110100100000", -- 7455 FREE #<CONS 0 7456>
 "00000000000000000001110100100001", -- 7456 FREE #<CONS 0 7457>
 "00000000000000000001110100100010", -- 7457 FREE #<CONS 0 7458>
 "00000000000000000001110100100011", -- 7458 FREE #<CONS 0 7459>
 "00000000000000000001110100100100", -- 7459 FREE #<CONS 0 7460>
 "00000000000000000001110100100101", -- 7460 FREE #<CONS 0 7461>
 "00000000000000000001110100100110", -- 7461 FREE #<CONS 0 7462>
 "00000000000000000001110100100111", -- 7462 FREE #<CONS 0 7463>
 "00000000000000000001110100101000", -- 7463 FREE #<CONS 0 7464>
 "00000000000000000001110100101001", -- 7464 FREE #<CONS 0 7465>
 "00000000000000000001110100101010", -- 7465 FREE #<CONS 0 7466>
 "00000000000000000001110100101011", -- 7466 FREE #<CONS 0 7467>
 "00000000000000000001110100101100", -- 7467 FREE #<CONS 0 7468>
 "00000000000000000001110100101101", -- 7468 FREE #<CONS 0 7469>
 "00000000000000000001110100101110", -- 7469 FREE #<CONS 0 7470>
 "00000000000000000001110100101111", -- 7470 FREE #<CONS 0 7471>
 "00000000000000000001110100110000", -- 7471 FREE #<CONS 0 7472>
 "00000000000000000001110100110001", -- 7472 FREE #<CONS 0 7473>
 "00000000000000000001110100110010", -- 7473 FREE #<CONS 0 7474>
 "00000000000000000001110100110011", -- 7474 FREE #<CONS 0 7475>
 "00000000000000000001110100110100", -- 7475 FREE #<CONS 0 7476>
 "00000000000000000001110100110101", -- 7476 FREE #<CONS 0 7477>
 "00000000000000000001110100110110", -- 7477 FREE #<CONS 0 7478>
 "00000000000000000001110100110111", -- 7478 FREE #<CONS 0 7479>
 "00000000000000000001110100111000", -- 7479 FREE #<CONS 0 7480>
 "00000000000000000001110100111001", -- 7480 FREE #<CONS 0 7481>
 "00000000000000000001110100111010", -- 7481 FREE #<CONS 0 7482>
 "00000000000000000001110100111011", -- 7482 FREE #<CONS 0 7483>
 "00000000000000000001110100111100", -- 7483 FREE #<CONS 0 7484>
 "00000000000000000001110100111101", -- 7484 FREE #<CONS 0 7485>
 "00000000000000000001110100111110", -- 7485 FREE #<CONS 0 7486>
 "00000000000000000001110100111111", -- 7486 FREE #<CONS 0 7487>
 "00000000000000000001110101000000", -- 7487 FREE #<CONS 0 7488>
 "00000000000000000001110101000001", -- 7488 FREE #<CONS 0 7489>
 "00000000000000000001110101000010", -- 7489 FREE #<CONS 0 7490>
 "00000000000000000001110101000011", -- 7490 FREE #<CONS 0 7491>
 "00000000000000000001110101000100", -- 7491 FREE #<CONS 0 7492>
 "00000000000000000001110101000101", -- 7492 FREE #<CONS 0 7493>
 "00000000000000000001110101000110", -- 7493 FREE #<CONS 0 7494>
 "00000000000000000001110101000111", -- 7494 FREE #<CONS 0 7495>
 "00000000000000000001110101001000", -- 7495 FREE #<CONS 0 7496>
 "00000000000000000001110101001001", -- 7496 FREE #<CONS 0 7497>
 "00000000000000000001110101001010", -- 7497 FREE #<CONS 0 7498>
 "00000000000000000001110101001011", -- 7498 FREE #<CONS 0 7499>
 "00000000000000000001110101001100", -- 7499 FREE #<CONS 0 7500>
 "00000000000000000001110101001101", -- 7500 FREE #<CONS 0 7501>
 "00000000000000000001110101001110", -- 7501 FREE #<CONS 0 7502>
 "00000000000000000001110101001111", -- 7502 FREE #<CONS 0 7503>
 "00000000000000000001110101010000", -- 7503 FREE #<CONS 0 7504>
 "00000000000000000001110101010001", -- 7504 FREE #<CONS 0 7505>
 "00000000000000000001110101010010", -- 7505 FREE #<CONS 0 7506>
 "00000000000000000001110101010011", -- 7506 FREE #<CONS 0 7507>
 "00000000000000000001110101010100", -- 7507 FREE #<CONS 0 7508>
 "00000000000000000001110101010101", -- 7508 FREE #<CONS 0 7509>
 "00000000000000000001110101010110", -- 7509 FREE #<CONS 0 7510>
 "00000000000000000001110101010111", -- 7510 FREE #<CONS 0 7511>
 "00000000000000000001110101011000", -- 7511 FREE #<CONS 0 7512>
 "00000000000000000001110101011001", -- 7512 FREE #<CONS 0 7513>
 "00000000000000000001110101011010", -- 7513 FREE #<CONS 0 7514>
 "00000000000000000001110101011011", -- 7514 FREE #<CONS 0 7515>
 "00000000000000000001110101011100", -- 7515 FREE #<CONS 0 7516>
 "00000000000000000001110101011101", -- 7516 FREE #<CONS 0 7517>
 "00000000000000000001110101011110", -- 7517 FREE #<CONS 0 7518>
 "00000000000000000001110101011111", -- 7518 FREE #<CONS 0 7519>
 "00000000000000000001110101100000", -- 7519 FREE #<CONS 0 7520>
 "00000000000000000001110101100001", -- 7520 FREE #<CONS 0 7521>
 "00000000000000000001110101100010", -- 7521 FREE #<CONS 0 7522>
 "00000000000000000001110101100011", -- 7522 FREE #<CONS 0 7523>
 "00000000000000000001110101100100", -- 7523 FREE #<CONS 0 7524>
 "00000000000000000001110101100101", -- 7524 FREE #<CONS 0 7525>
 "00000000000000000001110101100110", -- 7525 FREE #<CONS 0 7526>
 "00000000000000000001110101100111", -- 7526 FREE #<CONS 0 7527>
 "00000000000000000001110101101000", -- 7527 FREE #<CONS 0 7528>
 "00000000000000000001110101101001", -- 7528 FREE #<CONS 0 7529>
 "00000000000000000001110101101010", -- 7529 FREE #<CONS 0 7530>
 "00000000000000000001110101101011", -- 7530 FREE #<CONS 0 7531>
 "00000000000000000001110101101100", -- 7531 FREE #<CONS 0 7532>
 "00000000000000000001110101101101", -- 7532 FREE #<CONS 0 7533>
 "00000000000000000001110101101110", -- 7533 FREE #<CONS 0 7534>
 "00000000000000000001110101101111", -- 7534 FREE #<CONS 0 7535>
 "00000000000000000001110101110000", -- 7535 FREE #<CONS 0 7536>
 "00000000000000000001110101110001", -- 7536 FREE #<CONS 0 7537>
 "00000000000000000001110101110010", -- 7537 FREE #<CONS 0 7538>
 "00000000000000000001110101110011", -- 7538 FREE #<CONS 0 7539>
 "00000000000000000001110101110100", -- 7539 FREE #<CONS 0 7540>
 "00000000000000000001110101110101", -- 7540 FREE #<CONS 0 7541>
 "00000000000000000001110101110110", -- 7541 FREE #<CONS 0 7542>
 "00000000000000000001110101110111", -- 7542 FREE #<CONS 0 7543>
 "00000000000000000001110101111000", -- 7543 FREE #<CONS 0 7544>
 "00000000000000000001110101111001", -- 7544 FREE #<CONS 0 7545>
 "00000000000000000001110101111010", -- 7545 FREE #<CONS 0 7546>
 "00000000000000000001110101111011", -- 7546 FREE #<CONS 0 7547>
 "00000000000000000001110101111100", -- 7547 FREE #<CONS 0 7548>
 "00000000000000000001110101111101", -- 7548 FREE #<CONS 0 7549>
 "00000000000000000001110101111110", -- 7549 FREE #<CONS 0 7550>
 "00000000000000000001110101111111", -- 7550 FREE #<CONS 0 7551>
 "00000000000000000001110110000000", -- 7551 FREE #<CONS 0 7552>
 "00000000000000000001110110000001", -- 7552 FREE #<CONS 0 7553>
 "00000000000000000001110110000010", -- 7553 FREE #<CONS 0 7554>
 "00000000000000000001110110000011", -- 7554 FREE #<CONS 0 7555>
 "00000000000000000001110110000100", -- 7555 FREE #<CONS 0 7556>
 "00000000000000000001110110000101", -- 7556 FREE #<CONS 0 7557>
 "00000000000000000001110110000110", -- 7557 FREE #<CONS 0 7558>
 "00000000000000000001110110000111", -- 7558 FREE #<CONS 0 7559>
 "00000000000000000001110110001000", -- 7559 FREE #<CONS 0 7560>
 "00000000000000000001110110001001", -- 7560 FREE #<CONS 0 7561>
 "00000000000000000001110110001010", -- 7561 FREE #<CONS 0 7562>
 "00000000000000000001110110001011", -- 7562 FREE #<CONS 0 7563>
 "00000000000000000001110110001100", -- 7563 FREE #<CONS 0 7564>
 "00000000000000000001110110001101", -- 7564 FREE #<CONS 0 7565>
 "00000000000000000001110110001110", -- 7565 FREE #<CONS 0 7566>
 "00000000000000000001110110001111", -- 7566 FREE #<CONS 0 7567>
 "00000000000000000001110110010000", -- 7567 FREE #<CONS 0 7568>
 "00000000000000000001110110010001", -- 7568 FREE #<CONS 0 7569>
 "00000000000000000001110110010010", -- 7569 FREE #<CONS 0 7570>
 "00000000000000000001110110010011", -- 7570 FREE #<CONS 0 7571>
 "00000000000000000001110110010100", -- 7571 FREE #<CONS 0 7572>
 "00000000000000000001110110010101", -- 7572 FREE #<CONS 0 7573>
 "00000000000000000001110110010110", -- 7573 FREE #<CONS 0 7574>
 "00000000000000000001110110010111", -- 7574 FREE #<CONS 0 7575>
 "00000000000000000001110110011000", -- 7575 FREE #<CONS 0 7576>
 "00000000000000000001110110011001", -- 7576 FREE #<CONS 0 7577>
 "00000000000000000001110110011010", -- 7577 FREE #<CONS 0 7578>
 "00000000000000000001110110011011", -- 7578 FREE #<CONS 0 7579>
 "00000000000000000001110110011100", -- 7579 FREE #<CONS 0 7580>
 "00000000000000000001110110011101", -- 7580 FREE #<CONS 0 7581>
 "00000000000000000001110110011110", -- 7581 FREE #<CONS 0 7582>
 "00000000000000000001110110011111", -- 7582 FREE #<CONS 0 7583>
 "00000000000000000001110110100000", -- 7583 FREE #<CONS 0 7584>
 "00000000000000000001110110100001", -- 7584 FREE #<CONS 0 7585>
 "00000000000000000001110110100010", -- 7585 FREE #<CONS 0 7586>
 "00000000000000000001110110100011", -- 7586 FREE #<CONS 0 7587>
 "00000000000000000001110110100100", -- 7587 FREE #<CONS 0 7588>
 "00000000000000000001110110100101", -- 7588 FREE #<CONS 0 7589>
 "00000000000000000001110110100110", -- 7589 FREE #<CONS 0 7590>
 "00000000000000000001110110100111", -- 7590 FREE #<CONS 0 7591>
 "00000000000000000001110110101000", -- 7591 FREE #<CONS 0 7592>
 "00000000000000000001110110101001", -- 7592 FREE #<CONS 0 7593>
 "00000000000000000001110110101010", -- 7593 FREE #<CONS 0 7594>
 "00000000000000000001110110101011", -- 7594 FREE #<CONS 0 7595>
 "00000000000000000001110110101100", -- 7595 FREE #<CONS 0 7596>
 "00000000000000000001110110101101", -- 7596 FREE #<CONS 0 7597>
 "00000000000000000001110110101110", -- 7597 FREE #<CONS 0 7598>
 "00000000000000000001110110101111", -- 7598 FREE #<CONS 0 7599>
 "00000000000000000001110110110000", -- 7599 FREE #<CONS 0 7600>
 "00000000000000000001110110110001", -- 7600 FREE #<CONS 0 7601>
 "00000000000000000001110110110010", -- 7601 FREE #<CONS 0 7602>
 "00000000000000000001110110110011", -- 7602 FREE #<CONS 0 7603>
 "00000000000000000001110110110100", -- 7603 FREE #<CONS 0 7604>
 "00000000000000000001110110110101", -- 7604 FREE #<CONS 0 7605>
 "00000000000000000001110110110110", -- 7605 FREE #<CONS 0 7606>
 "00000000000000000001110110110111", -- 7606 FREE #<CONS 0 7607>
 "00000000000000000001110110111000", -- 7607 FREE #<CONS 0 7608>
 "00000000000000000001110110111001", -- 7608 FREE #<CONS 0 7609>
 "00000000000000000001110110111010", -- 7609 FREE #<CONS 0 7610>
 "00000000000000000001110110111011", -- 7610 FREE #<CONS 0 7611>
 "00000000000000000001110110111100", -- 7611 FREE #<CONS 0 7612>
 "00000000000000000001110110111101", -- 7612 FREE #<CONS 0 7613>
 "00000000000000000001110110111110", -- 7613 FREE #<CONS 0 7614>
 "00000000000000000001110110111111", -- 7614 FREE #<CONS 0 7615>
 "00000000000000000001110111000000", -- 7615 FREE #<CONS 0 7616>
 "00000000000000000001110111000001", -- 7616 FREE #<CONS 0 7617>
 "00000000000000000001110111000010", -- 7617 FREE #<CONS 0 7618>
 "00000000000000000001110111000011", -- 7618 FREE #<CONS 0 7619>
 "00000000000000000001110111000100", -- 7619 FREE #<CONS 0 7620>
 "00000000000000000001110111000101", -- 7620 FREE #<CONS 0 7621>
 "00000000000000000001110111000110", -- 7621 FREE #<CONS 0 7622>
 "00000000000000000001110111000111", -- 7622 FREE #<CONS 0 7623>
 "00000000000000000001110111001000", -- 7623 FREE #<CONS 0 7624>
 "00000000000000000001110111001001", -- 7624 FREE #<CONS 0 7625>
 "00000000000000000001110111001010", -- 7625 FREE #<CONS 0 7626>
 "00000000000000000001110111001011", -- 7626 FREE #<CONS 0 7627>
 "00000000000000000001110111001100", -- 7627 FREE #<CONS 0 7628>
 "00000000000000000001110111001101", -- 7628 FREE #<CONS 0 7629>
 "00000000000000000001110111001110", -- 7629 FREE #<CONS 0 7630>
 "00000000000000000001110111001111", -- 7630 FREE #<CONS 0 7631>
 "00000000000000000001110111010000", -- 7631 FREE #<CONS 0 7632>
 "00000000000000000001110111010001", -- 7632 FREE #<CONS 0 7633>
 "00000000000000000001110111010010", -- 7633 FREE #<CONS 0 7634>
 "00000000000000000001110111010011", -- 7634 FREE #<CONS 0 7635>
 "00000000000000000001110111010100", -- 7635 FREE #<CONS 0 7636>
 "00000000000000000001110111010101", -- 7636 FREE #<CONS 0 7637>
 "00000000000000000001110111010110", -- 7637 FREE #<CONS 0 7638>
 "00000000000000000001110111010111", -- 7638 FREE #<CONS 0 7639>
 "00000000000000000001110111011000", -- 7639 FREE #<CONS 0 7640>
 "00000000000000000001110111011001", -- 7640 FREE #<CONS 0 7641>
 "00000000000000000001110111011010", -- 7641 FREE #<CONS 0 7642>
 "00000000000000000001110111011011", -- 7642 FREE #<CONS 0 7643>
 "00000000000000000001110111011100", -- 7643 FREE #<CONS 0 7644>
 "00000000000000000001110111011101", -- 7644 FREE #<CONS 0 7645>
 "00000000000000000001110111011110", -- 7645 FREE #<CONS 0 7646>
 "00000000000000000001110111011111", -- 7646 FREE #<CONS 0 7647>
 "00000000000000000001110111100000", -- 7647 FREE #<CONS 0 7648>
 "00000000000000000001110111100001", -- 7648 FREE #<CONS 0 7649>
 "00000000000000000001110111100010", -- 7649 FREE #<CONS 0 7650>
 "00000000000000000001110111100011", -- 7650 FREE #<CONS 0 7651>
 "00000000000000000001110111100100", -- 7651 FREE #<CONS 0 7652>
 "00000000000000000001110111100101", -- 7652 FREE #<CONS 0 7653>
 "00000000000000000001110111100110", -- 7653 FREE #<CONS 0 7654>
 "00000000000000000001110111100111", -- 7654 FREE #<CONS 0 7655>
 "00000000000000000001110111101000", -- 7655 FREE #<CONS 0 7656>
 "00000000000000000001110111101001", -- 7656 FREE #<CONS 0 7657>
 "00000000000000000001110111101010", -- 7657 FREE #<CONS 0 7658>
 "00000000000000000001110111101011", -- 7658 FREE #<CONS 0 7659>
 "00000000000000000001110111101100", -- 7659 FREE #<CONS 0 7660>
 "00000000000000000001110111101101", -- 7660 FREE #<CONS 0 7661>
 "00000000000000000001110111101110", -- 7661 FREE #<CONS 0 7662>
 "00000000000000000001110111101111", -- 7662 FREE #<CONS 0 7663>
 "00000000000000000001110111110000", -- 7663 FREE #<CONS 0 7664>
 "00000000000000000001110111110001", -- 7664 FREE #<CONS 0 7665>
 "00000000000000000001110111110010", -- 7665 FREE #<CONS 0 7666>
 "00000000000000000001110111110011", -- 7666 FREE #<CONS 0 7667>
 "00000000000000000001110111110100", -- 7667 FREE #<CONS 0 7668>
 "00000000000000000001110111110101", -- 7668 FREE #<CONS 0 7669>
 "00000000000000000001110111110110", -- 7669 FREE #<CONS 0 7670>
 "00000000000000000001110111110111", -- 7670 FREE #<CONS 0 7671>
 "00000000000000000001110111111000", -- 7671 FREE #<CONS 0 7672>
 "00000000000000000001110111111001", -- 7672 FREE #<CONS 0 7673>
 "00000000000000000001110111111010", -- 7673 FREE #<CONS 0 7674>
 "00000000000000000001110111111011", -- 7674 FREE #<CONS 0 7675>
 "00000000000000000001110111111100", -- 7675 FREE #<CONS 0 7676>
 "00000000000000000001110111111101", -- 7676 FREE #<CONS 0 7677>
 "00000000000000000001110111111110", -- 7677 FREE #<CONS 0 7678>
 "00000000000000000001110111111111", -- 7678 FREE #<CONS 0 7679>
 "00000000000000000001111000000000", -- 7679 FREE #<CONS 0 7680>
 "00000000000000000001111000000001", -- 7680 FREE #<CONS 0 7681>
 "00000000000000000001111000000010", -- 7681 FREE #<CONS 0 7682>
 "00000000000000000001111000000011", -- 7682 FREE #<CONS 0 7683>
 "00000000000000000001111000000100", -- 7683 FREE #<CONS 0 7684>
 "00000000000000000001111000000101", -- 7684 FREE #<CONS 0 7685>
 "00000000000000000001111000000110", -- 7685 FREE #<CONS 0 7686>
 "00000000000000000001111000000111", -- 7686 FREE #<CONS 0 7687>
 "00000000000000000001111000001000", -- 7687 FREE #<CONS 0 7688>
 "00000000000000000001111000001001", -- 7688 FREE #<CONS 0 7689>
 "00000000000000000001111000001010", -- 7689 FREE #<CONS 0 7690>
 "00000000000000000001111000001011", -- 7690 FREE #<CONS 0 7691>
 "00000000000000000001111000001100", -- 7691 FREE #<CONS 0 7692>
 "00000000000000000001111000001101", -- 7692 FREE #<CONS 0 7693>
 "00000000000000000001111000001110", -- 7693 FREE #<CONS 0 7694>
 "00000000000000000001111000001111", -- 7694 FREE #<CONS 0 7695>
 "00000000000000000001111000010000", -- 7695 FREE #<CONS 0 7696>
 "00000000000000000001111000010001", -- 7696 FREE #<CONS 0 7697>
 "00000000000000000001111000010010", -- 7697 FREE #<CONS 0 7698>
 "00000000000000000001111000010011", -- 7698 FREE #<CONS 0 7699>
 "00000000000000000001111000010100", -- 7699 FREE #<CONS 0 7700>
 "00000000000000000001111000010101", -- 7700 FREE #<CONS 0 7701>
 "00000000000000000001111000010110", -- 7701 FREE #<CONS 0 7702>
 "00000000000000000001111000010111", -- 7702 FREE #<CONS 0 7703>
 "00000000000000000001111000011000", -- 7703 FREE #<CONS 0 7704>
 "00000000000000000001111000011001", -- 7704 FREE #<CONS 0 7705>
 "00000000000000000001111000011010", -- 7705 FREE #<CONS 0 7706>
 "00000000000000000001111000011011", -- 7706 FREE #<CONS 0 7707>
 "00000000000000000001111000011100", -- 7707 FREE #<CONS 0 7708>
 "00000000000000000001111000011101", -- 7708 FREE #<CONS 0 7709>
 "00000000000000000001111000011110", -- 7709 FREE #<CONS 0 7710>
 "00000000000000000001111000011111", -- 7710 FREE #<CONS 0 7711>
 "00000000000000000001111000100000", -- 7711 FREE #<CONS 0 7712>
 "00000000000000000001111000100001", -- 7712 FREE #<CONS 0 7713>
 "00000000000000000001111000100010", -- 7713 FREE #<CONS 0 7714>
 "00000000000000000001111000100011", -- 7714 FREE #<CONS 0 7715>
 "00000000000000000001111000100100", -- 7715 FREE #<CONS 0 7716>
 "00000000000000000001111000100101", -- 7716 FREE #<CONS 0 7717>
 "00000000000000000001111000100110", -- 7717 FREE #<CONS 0 7718>
 "00000000000000000001111000100111", -- 7718 FREE #<CONS 0 7719>
 "00000000000000000001111000101000", -- 7719 FREE #<CONS 0 7720>
 "00000000000000000001111000101001", -- 7720 FREE #<CONS 0 7721>
 "00000000000000000001111000101010", -- 7721 FREE #<CONS 0 7722>
 "00000000000000000001111000101011", -- 7722 FREE #<CONS 0 7723>
 "00000000000000000001111000101100", -- 7723 FREE #<CONS 0 7724>
 "00000000000000000001111000101101", -- 7724 FREE #<CONS 0 7725>
 "00000000000000000001111000101110", -- 7725 FREE #<CONS 0 7726>
 "00000000000000000001111000101111", -- 7726 FREE #<CONS 0 7727>
 "00000000000000000001111000110000", -- 7727 FREE #<CONS 0 7728>
 "00000000000000000001111000110001", -- 7728 FREE #<CONS 0 7729>
 "00000000000000000001111000110010", -- 7729 FREE #<CONS 0 7730>
 "00000000000000000001111000110011", -- 7730 FREE #<CONS 0 7731>
 "00000000000000000001111000110100", -- 7731 FREE #<CONS 0 7732>
 "00000000000000000001111000110101", -- 7732 FREE #<CONS 0 7733>
 "00000000000000000001111000110110", -- 7733 FREE #<CONS 0 7734>
 "00000000000000000001111000110111", -- 7734 FREE #<CONS 0 7735>
 "00000000000000000001111000111000", -- 7735 FREE #<CONS 0 7736>
 "00000000000000000001111000111001", -- 7736 FREE #<CONS 0 7737>
 "00000000000000000001111000111010", -- 7737 FREE #<CONS 0 7738>
 "00000000000000000001111000111011", -- 7738 FREE #<CONS 0 7739>
 "00000000000000000001111000111100", -- 7739 FREE #<CONS 0 7740>
 "00000000000000000001111000111101", -- 7740 FREE #<CONS 0 7741>
 "00000000000000000001111000111110", -- 7741 FREE #<CONS 0 7742>
 "00000000000000000001111000111111", -- 7742 FREE #<CONS 0 7743>
 "00000000000000000001111001000000", -- 7743 FREE #<CONS 0 7744>
 "00000000000000000001111001000001", -- 7744 FREE #<CONS 0 7745>
 "00000000000000000001111001000010", -- 7745 FREE #<CONS 0 7746>
 "00000000000000000001111001000011", -- 7746 FREE #<CONS 0 7747>
 "00000000000000000001111001000100", -- 7747 FREE #<CONS 0 7748>
 "00000000000000000001111001000101", -- 7748 FREE #<CONS 0 7749>
 "00000000000000000001111001000110", -- 7749 FREE #<CONS 0 7750>
 "00000000000000000001111001000111", -- 7750 FREE #<CONS 0 7751>
 "00000000000000000001111001001000", -- 7751 FREE #<CONS 0 7752>
 "00000000000000000001111001001001", -- 7752 FREE #<CONS 0 7753>
 "00000000000000000001111001001010", -- 7753 FREE #<CONS 0 7754>
 "00000000000000000001111001001011", -- 7754 FREE #<CONS 0 7755>
 "00000000000000000001111001001100", -- 7755 FREE #<CONS 0 7756>
 "00000000000000000001111001001101", -- 7756 FREE #<CONS 0 7757>
 "00000000000000000001111001001110", -- 7757 FREE #<CONS 0 7758>
 "00000000000000000001111001001111", -- 7758 FREE #<CONS 0 7759>
 "00000000000000000001111001010000", -- 7759 FREE #<CONS 0 7760>
 "00000000000000000001111001010001", -- 7760 FREE #<CONS 0 7761>
 "00000000000000000001111001010010", -- 7761 FREE #<CONS 0 7762>
 "00000000000000000001111001010011", -- 7762 FREE #<CONS 0 7763>
 "00000000000000000001111001010100", -- 7763 FREE #<CONS 0 7764>
 "00000000000000000001111001010101", -- 7764 FREE #<CONS 0 7765>
 "00000000000000000001111001010110", -- 7765 FREE #<CONS 0 7766>
 "00000000000000000001111001010111", -- 7766 FREE #<CONS 0 7767>
 "00000000000000000001111001011000", -- 7767 FREE #<CONS 0 7768>
 "00000000000000000001111001011001", -- 7768 FREE #<CONS 0 7769>
 "00000000000000000001111001011010", -- 7769 FREE #<CONS 0 7770>
 "00000000000000000001111001011011", -- 7770 FREE #<CONS 0 7771>
 "00000000000000000001111001011100", -- 7771 FREE #<CONS 0 7772>
 "00000000000000000001111001011101", -- 7772 FREE #<CONS 0 7773>
 "00000000000000000001111001011110", -- 7773 FREE #<CONS 0 7774>
 "00000000000000000001111001011111", -- 7774 FREE #<CONS 0 7775>
 "00000000000000000001111001100000", -- 7775 FREE #<CONS 0 7776>
 "00000000000000000001111001100001", -- 7776 FREE #<CONS 0 7777>
 "00000000000000000001111001100010", -- 7777 FREE #<CONS 0 7778>
 "00000000000000000001111001100011", -- 7778 FREE #<CONS 0 7779>
 "00000000000000000001111001100100", -- 7779 FREE #<CONS 0 7780>
 "00000000000000000001111001100101", -- 7780 FREE #<CONS 0 7781>
 "00000000000000000001111001100110", -- 7781 FREE #<CONS 0 7782>
 "00000000000000000001111001100111", -- 7782 FREE #<CONS 0 7783>
 "00000000000000000001111001101000", -- 7783 FREE #<CONS 0 7784>
 "00000000000000000001111001101001", -- 7784 FREE #<CONS 0 7785>
 "00000000000000000001111001101010", -- 7785 FREE #<CONS 0 7786>
 "00000000000000000001111001101011", -- 7786 FREE #<CONS 0 7787>
 "00000000000000000001111001101100", -- 7787 FREE #<CONS 0 7788>
 "00000000000000000001111001101101", -- 7788 FREE #<CONS 0 7789>
 "00000000000000000001111001101110", -- 7789 FREE #<CONS 0 7790>
 "00000000000000000001111001101111", -- 7790 FREE #<CONS 0 7791>
 "00000000000000000001111001110000", -- 7791 FREE #<CONS 0 7792>
 "00000000000000000001111001110001", -- 7792 FREE #<CONS 0 7793>
 "00000000000000000001111001110010", -- 7793 FREE #<CONS 0 7794>
 "00000000000000000001111001110011", -- 7794 FREE #<CONS 0 7795>
 "00000000000000000001111001110100", -- 7795 FREE #<CONS 0 7796>
 "00000000000000000001111001110101", -- 7796 FREE #<CONS 0 7797>
 "00000000000000000001111001110110", -- 7797 FREE #<CONS 0 7798>
 "00000000000000000001111001110111", -- 7798 FREE #<CONS 0 7799>
 "00000000000000000001111001111000", -- 7799 FREE #<CONS 0 7800>
 "00000000000000000001111001111001", -- 7800 FREE #<CONS 0 7801>
 "00000000000000000001111001111010", -- 7801 FREE #<CONS 0 7802>
 "00000000000000000001111001111011", -- 7802 FREE #<CONS 0 7803>
 "00000000000000000001111001111100", -- 7803 FREE #<CONS 0 7804>
 "00000000000000000001111001111101", -- 7804 FREE #<CONS 0 7805>
 "00000000000000000001111001111110", -- 7805 FREE #<CONS 0 7806>
 "00000000000000000001111001111111", -- 7806 FREE #<CONS 0 7807>
 "00000000000000000001111010000000", -- 7807 FREE #<CONS 0 7808>
 "00000000000000000001111010000001", -- 7808 FREE #<CONS 0 7809>
 "00000000000000000001111010000010", -- 7809 FREE #<CONS 0 7810>
 "00000000000000000001111010000011", -- 7810 FREE #<CONS 0 7811>
 "00000000000000000001111010000100", -- 7811 FREE #<CONS 0 7812>
 "00000000000000000001111010000101", -- 7812 FREE #<CONS 0 7813>
 "00000000000000000001111010000110", -- 7813 FREE #<CONS 0 7814>
 "00000000000000000001111010000111", -- 7814 FREE #<CONS 0 7815>
 "00000000000000000001111010001000", -- 7815 FREE #<CONS 0 7816>
 "00000000000000000001111010001001", -- 7816 FREE #<CONS 0 7817>
 "00000000000000000001111010001010", -- 7817 FREE #<CONS 0 7818>
 "00000000000000000001111010001011", -- 7818 FREE #<CONS 0 7819>
 "00000000000000000001111010001100", -- 7819 FREE #<CONS 0 7820>
 "00000000000000000001111010001101", -- 7820 FREE #<CONS 0 7821>
 "00000000000000000001111010001110", -- 7821 FREE #<CONS 0 7822>
 "00000000000000000001111010001111", -- 7822 FREE #<CONS 0 7823>
 "00000000000000000001111010010000", -- 7823 FREE #<CONS 0 7824>
 "00000000000000000001111010010001", -- 7824 FREE #<CONS 0 7825>
 "00000000000000000001111010010010", -- 7825 FREE #<CONS 0 7826>
 "00000000000000000001111010010011", -- 7826 FREE #<CONS 0 7827>
 "00000000000000000001111010010100", -- 7827 FREE #<CONS 0 7828>
 "00000000000000000001111010010101", -- 7828 FREE #<CONS 0 7829>
 "00000000000000000001111010010110", -- 7829 FREE #<CONS 0 7830>
 "00000000000000000001111010010111", -- 7830 FREE #<CONS 0 7831>
 "00000000000000000001111010011000", -- 7831 FREE #<CONS 0 7832>
 "00000000000000000001111010011001", -- 7832 FREE #<CONS 0 7833>
 "00000000000000000001111010011010", -- 7833 FREE #<CONS 0 7834>
 "00000000000000000001111010011011", -- 7834 FREE #<CONS 0 7835>
 "00000000000000000001111010011100", -- 7835 FREE #<CONS 0 7836>
 "00000000000000000001111010011101", -- 7836 FREE #<CONS 0 7837>
 "00000000000000000001111010011110", -- 7837 FREE #<CONS 0 7838>
 "00000000000000000001111010011111", -- 7838 FREE #<CONS 0 7839>
 "00000000000000000001111010100000", -- 7839 FREE #<CONS 0 7840>
 "00000000000000000001111010100001", -- 7840 FREE #<CONS 0 7841>
 "00000000000000000001111010100010", -- 7841 FREE #<CONS 0 7842>
 "00000000000000000001111010100011", -- 7842 FREE #<CONS 0 7843>
 "00000000000000000001111010100100", -- 7843 FREE #<CONS 0 7844>
 "00000000000000000001111010100101", -- 7844 FREE #<CONS 0 7845>
 "00000000000000000001111010100110", -- 7845 FREE #<CONS 0 7846>
 "00000000000000000001111010100111", -- 7846 FREE #<CONS 0 7847>
 "00000000000000000001111010101000", -- 7847 FREE #<CONS 0 7848>
 "00000000000000000001111010101001", -- 7848 FREE #<CONS 0 7849>
 "00000000000000000001111010101010", -- 7849 FREE #<CONS 0 7850>
 "00000000000000000001111010101011", -- 7850 FREE #<CONS 0 7851>
 "00000000000000000001111010101100", -- 7851 FREE #<CONS 0 7852>
 "00000000000000000001111010101101", -- 7852 FREE #<CONS 0 7853>
 "00000000000000000001111010101110", -- 7853 FREE #<CONS 0 7854>
 "00000000000000000001111010101111", -- 7854 FREE #<CONS 0 7855>
 "00000000000000000001111010110000", -- 7855 FREE #<CONS 0 7856>
 "00000000000000000001111010110001", -- 7856 FREE #<CONS 0 7857>
 "00000000000000000001111010110010", -- 7857 FREE #<CONS 0 7858>
 "00000000000000000001111010110011", -- 7858 FREE #<CONS 0 7859>
 "00000000000000000001111010110100", -- 7859 FREE #<CONS 0 7860>
 "00000000000000000001111010110101", -- 7860 FREE #<CONS 0 7861>
 "00000000000000000001111010110110", -- 7861 FREE #<CONS 0 7862>
 "00000000000000000001111010110111", -- 7862 FREE #<CONS 0 7863>
 "00000000000000000001111010111000", -- 7863 FREE #<CONS 0 7864>
 "00000000000000000001111010111001", -- 7864 FREE #<CONS 0 7865>
 "00000000000000000001111010111010", -- 7865 FREE #<CONS 0 7866>
 "00000000000000000001111010111011", -- 7866 FREE #<CONS 0 7867>
 "00000000000000000001111010111100", -- 7867 FREE #<CONS 0 7868>
 "00000000000000000001111010111101", -- 7868 FREE #<CONS 0 7869>
 "00000000000000000001111010111110", -- 7869 FREE #<CONS 0 7870>
 "00000000000000000001111010111111", -- 7870 FREE #<CONS 0 7871>
 "00000000000000000001111011000000", -- 7871 FREE #<CONS 0 7872>
 "00000000000000000001111011000001", -- 7872 FREE #<CONS 0 7873>
 "00000000000000000001111011000010", -- 7873 FREE #<CONS 0 7874>
 "00000000000000000001111011000011", -- 7874 FREE #<CONS 0 7875>
 "00000000000000000001111011000100", -- 7875 FREE #<CONS 0 7876>
 "00000000000000000001111011000101", -- 7876 FREE #<CONS 0 7877>
 "00000000000000000001111011000110", -- 7877 FREE #<CONS 0 7878>
 "00000000000000000001111011000111", -- 7878 FREE #<CONS 0 7879>
 "00000000000000000001111011001000", -- 7879 FREE #<CONS 0 7880>
 "00000000000000000001111011001001", -- 7880 FREE #<CONS 0 7881>
 "00000000000000000001111011001010", -- 7881 FREE #<CONS 0 7882>
 "00000000000000000001111011001011", -- 7882 FREE #<CONS 0 7883>
 "00000000000000000001111011001100", -- 7883 FREE #<CONS 0 7884>
 "00000000000000000001111011001101", -- 7884 FREE #<CONS 0 7885>
 "00000000000000000001111011001110", -- 7885 FREE #<CONS 0 7886>
 "00000000000000000001111011001111", -- 7886 FREE #<CONS 0 7887>
 "00000000000000000001111011010000", -- 7887 FREE #<CONS 0 7888>
 "00000000000000000001111011010001", -- 7888 FREE #<CONS 0 7889>
 "00000000000000000001111011010010", -- 7889 FREE #<CONS 0 7890>
 "00000000000000000001111011010011", -- 7890 FREE #<CONS 0 7891>
 "00000000000000000001111011010100", -- 7891 FREE #<CONS 0 7892>
 "00000000000000000001111011010101", -- 7892 FREE #<CONS 0 7893>
 "00000000000000000001111011010110", -- 7893 FREE #<CONS 0 7894>
 "00000000000000000001111011010111", -- 7894 FREE #<CONS 0 7895>
 "00000000000000000001111011011000", -- 7895 FREE #<CONS 0 7896>
 "00000000000000000001111011011001", -- 7896 FREE #<CONS 0 7897>
 "00000000000000000001111011011010", -- 7897 FREE #<CONS 0 7898>
 "00000000000000000001111011011011", -- 7898 FREE #<CONS 0 7899>
 "00000000000000000001111011011100", -- 7899 FREE #<CONS 0 7900>
 "00000000000000000001111011011101", -- 7900 FREE #<CONS 0 7901>
 "00000000000000000001111011011110", -- 7901 FREE #<CONS 0 7902>
 "00000000000000000001111011011111", -- 7902 FREE #<CONS 0 7903>
 "00000000000000000001111011100000", -- 7903 FREE #<CONS 0 7904>
 "00000000000000000001111011100001", -- 7904 FREE #<CONS 0 7905>
 "00000000000000000001111011100010", -- 7905 FREE #<CONS 0 7906>
 "00000000000000000001111011100011", -- 7906 FREE #<CONS 0 7907>
 "00000000000000000001111011100100", -- 7907 FREE #<CONS 0 7908>
 "00000000000000000001111011100101", -- 7908 FREE #<CONS 0 7909>
 "00000000000000000001111011100110", -- 7909 FREE #<CONS 0 7910>
 "00000000000000000001111011100111", -- 7910 FREE #<CONS 0 7911>
 "00000000000000000001111011101000", -- 7911 FREE #<CONS 0 7912>
 "00000000000000000001111011101001", -- 7912 FREE #<CONS 0 7913>
 "00000000000000000001111011101010", -- 7913 FREE #<CONS 0 7914>
 "00000000000000000001111011101011", -- 7914 FREE #<CONS 0 7915>
 "00000000000000000001111011101100", -- 7915 FREE #<CONS 0 7916>
 "00000000000000000001111011101101", -- 7916 FREE #<CONS 0 7917>
 "00000000000000000001111011101110", -- 7917 FREE #<CONS 0 7918>
 "00000000000000000001111011101111", -- 7918 FREE #<CONS 0 7919>
 "00000000000000000001111011110000", -- 7919 FREE #<CONS 0 7920>
 "00000000000000000001111011110001", -- 7920 FREE #<CONS 0 7921>
 "00000000000000000001111011110010", -- 7921 FREE #<CONS 0 7922>
 "00000000000000000001111011110011", -- 7922 FREE #<CONS 0 7923>
 "00000000000000000001111011110100", -- 7923 FREE #<CONS 0 7924>
 "00000000000000000001111011110101", -- 7924 FREE #<CONS 0 7925>
 "00000000000000000001111011110110", -- 7925 FREE #<CONS 0 7926>
 "00000000000000000001111011110111", -- 7926 FREE #<CONS 0 7927>
 "00000000000000000001111011111000", -- 7927 FREE #<CONS 0 7928>
 "00000000000000000001111011111001", -- 7928 FREE #<CONS 0 7929>
 "00000000000000000001111011111010", -- 7929 FREE #<CONS 0 7930>
 "00000000000000000001111011111011", -- 7930 FREE #<CONS 0 7931>
 "00000000000000000001111011111100", -- 7931 FREE #<CONS 0 7932>
 "00000000000000000001111011111101", -- 7932 FREE #<CONS 0 7933>
 "00000000000000000001111011111110", -- 7933 FREE #<CONS 0 7934>
 "00000000000000000001111011111111", -- 7934 FREE #<CONS 0 7935>
 "00000000000000000001111100000000", -- 7935 FREE #<CONS 0 7936>
 "00000000000000000001111100000001", -- 7936 FREE #<CONS 0 7937>
 "00000000000000000001111100000010", -- 7937 FREE #<CONS 0 7938>
 "00000000000000000001111100000011", -- 7938 FREE #<CONS 0 7939>
 "00000000000000000001111100000100", -- 7939 FREE #<CONS 0 7940>
 "00000000000000000001111100000101", -- 7940 FREE #<CONS 0 7941>
 "00000000000000000001111100000110", -- 7941 FREE #<CONS 0 7942>
 "00000000000000000001111100000111", -- 7942 FREE #<CONS 0 7943>
 "00000000000000000001111100001000", -- 7943 FREE #<CONS 0 7944>
 "00000000000000000001111100001001", -- 7944 FREE #<CONS 0 7945>
 "00000000000000000001111100001010", -- 7945 FREE #<CONS 0 7946>
 "00000000000000000001111100001011", -- 7946 FREE #<CONS 0 7947>
 "00000000000000000001111100001100", -- 7947 FREE #<CONS 0 7948>
 "00000000000000000001111100001101", -- 7948 FREE #<CONS 0 7949>
 "00000000000000000001111100001110", -- 7949 FREE #<CONS 0 7950>
 "00000000000000000001111100001111", -- 7950 FREE #<CONS 0 7951>
 "00000000000000000001111100010000", -- 7951 FREE #<CONS 0 7952>
 "00000000000000000001111100010001", -- 7952 FREE #<CONS 0 7953>
 "00000000000000000001111100010010", -- 7953 FREE #<CONS 0 7954>
 "00000000000000000001111100010011", -- 7954 FREE #<CONS 0 7955>
 "00000000000000000001111100010100", -- 7955 FREE #<CONS 0 7956>
 "00000000000000000001111100010101", -- 7956 FREE #<CONS 0 7957>
 "00000000000000000001111100010110", -- 7957 FREE #<CONS 0 7958>
 "00000000000000000001111100010111", -- 7958 FREE #<CONS 0 7959>
 "00000000000000000001111100011000", -- 7959 FREE #<CONS 0 7960>
 "00000000000000000001111100011001", -- 7960 FREE #<CONS 0 7961>
 "00000000000000000001111100011010", -- 7961 FREE #<CONS 0 7962>
 "00000000000000000001111100011011", -- 7962 FREE #<CONS 0 7963>
 "00000000000000000001111100011100", -- 7963 FREE #<CONS 0 7964>
 "00000000000000000001111100011101", -- 7964 FREE #<CONS 0 7965>
 "00000000000000000001111100011110", -- 7965 FREE #<CONS 0 7966>
 "00000000000000000001111100011111", -- 7966 FREE #<CONS 0 7967>
 "00000000000000000001111100100000", -- 7967 FREE #<CONS 0 7968>
 "00000000000000000001111100100001", -- 7968 FREE #<CONS 0 7969>
 "00000000000000000001111100100010", -- 7969 FREE #<CONS 0 7970>
 "00000000000000000001111100100011", -- 7970 FREE #<CONS 0 7971>
 "00000000000000000001111100100100", -- 7971 FREE #<CONS 0 7972>
 "00000000000000000001111100100101", -- 7972 FREE #<CONS 0 7973>
 "00000000000000000001111100100110", -- 7973 FREE #<CONS 0 7974>
 "00000000000000000001111100100111", -- 7974 FREE #<CONS 0 7975>
 "00000000000000000001111100101000", -- 7975 FREE #<CONS 0 7976>
 "00000000000000000001111100101001", -- 7976 FREE #<CONS 0 7977>
 "00000000000000000001111100101010", -- 7977 FREE #<CONS 0 7978>
 "00000000000000000001111100101011", -- 7978 FREE #<CONS 0 7979>
 "00000000000000000001111100101100", -- 7979 FREE #<CONS 0 7980>
 "00000000000000000001111100101101", -- 7980 FREE #<CONS 0 7981>
 "00000000000000000001111100101110", -- 7981 FREE #<CONS 0 7982>
 "00000000000000000001111100101111", -- 7982 FREE #<CONS 0 7983>
 "00000000000000000001111100110000", -- 7983 FREE #<CONS 0 7984>
 "00000000000000000001111100110001", -- 7984 FREE #<CONS 0 7985>
 "00000000000000000001111100110010", -- 7985 FREE #<CONS 0 7986>
 "00000000000000000001111100110011", -- 7986 FREE #<CONS 0 7987>
 "00000000000000000001111100110100", -- 7987 FREE #<CONS 0 7988>
 "00000000000000000001111100110101", -- 7988 FREE #<CONS 0 7989>
 "00000000000000000001111100110110", -- 7989 FREE #<CONS 0 7990>
 "00000000000000000001111100110111", -- 7990 FREE #<CONS 0 7991>
 "00000000000000000001111100111000", -- 7991 FREE #<CONS 0 7992>
 "00000000000000000001111100111001", -- 7992 FREE #<CONS 0 7993>
 "00000000000000000001111100111010", -- 7993 FREE #<CONS 0 7994>
 "00000000000000000001111100111011", -- 7994 FREE #<CONS 0 7995>
 "00000000000000000001111100111100", -- 7995 FREE #<CONS 0 7996>
 "00000000000000000001111100111101", -- 7996 FREE #<CONS 0 7997>
 "00000000000000000001111100111110", -- 7997 FREE #<CONS 0 7998>
 "00000000000000000001111100111111", -- 7998 FREE #<CONS 0 7999>
 "00000000000000000001111101000000", -- 7999 FREE #<CONS 0 8000>
 "00000000000000000001111101000001", -- 8000 FREE #<CONS 0 8001>
 "00000000000000000001111101000010", -- 8001 FREE #<CONS 0 8002>
 "00000000000000000001111101000011", -- 8002 FREE #<CONS 0 8003>
 "00000000000000000001111101000100", -- 8003 FREE #<CONS 0 8004>
 "00000000000000000001111101000101", -- 8004 FREE #<CONS 0 8005>
 "00000000000000000001111101000110", -- 8005 FREE #<CONS 0 8006>
 "00000000000000000001111101000111", -- 8006 FREE #<CONS 0 8007>
 "00000000000000000001111101001000", -- 8007 FREE #<CONS 0 8008>
 "00000000000000000001111101001001", -- 8008 FREE #<CONS 0 8009>
 "00000000000000000001111101001010", -- 8009 FREE #<CONS 0 8010>
 "00000000000000000001111101001011", -- 8010 FREE #<CONS 0 8011>
 "00000000000000000001111101001100", -- 8011 FREE #<CONS 0 8012>
 "00000000000000000001111101001101", -- 8012 FREE #<CONS 0 8013>
 "00000000000000000001111101001110", -- 8013 FREE #<CONS 0 8014>
 "00000000000000000001111101001111", -- 8014 FREE #<CONS 0 8015>
 "00000000000000000001111101010000", -- 8015 FREE #<CONS 0 8016>
 "00000000000000000001111101010001", -- 8016 FREE #<CONS 0 8017>
 "00000000000000000001111101010010", -- 8017 FREE #<CONS 0 8018>
 "00000000000000000001111101010011", -- 8018 FREE #<CONS 0 8019>
 "00000000000000000001111101010100", -- 8019 FREE #<CONS 0 8020>
 "00000000000000000001111101010101", -- 8020 FREE #<CONS 0 8021>
 "00000000000000000001111101010110", -- 8021 FREE #<CONS 0 8022>
 "00000000000000000001111101010111", -- 8022 FREE #<CONS 0 8023>
 "00000000000000000001111101011000", -- 8023 FREE #<CONS 0 8024>
 "00000000000000000001111101011001", -- 8024 FREE #<CONS 0 8025>
 "00000000000000000001111101011010", -- 8025 FREE #<CONS 0 8026>
 "00000000000000000001111101011011", -- 8026 FREE #<CONS 0 8027>
 "00000000000000000001111101011100", -- 8027 FREE #<CONS 0 8028>
 "00000000000000000001111101011101", -- 8028 FREE #<CONS 0 8029>
 "00000000000000000001111101011110", -- 8029 FREE #<CONS 0 8030>
 "00000000000000000001111101011111", -- 8030 FREE #<CONS 0 8031>
 "00000000000000000001111101100000", -- 8031 FREE #<CONS 0 8032>
 "00000000000000000001111101100001", -- 8032 FREE #<CONS 0 8033>
 "00000000000000000001111101100010", -- 8033 FREE #<CONS 0 8034>
 "00000000000000000001111101100011", -- 8034 FREE #<CONS 0 8035>
 "00000000000000000001111101100100", -- 8035 FREE #<CONS 0 8036>
 "00000000000000000001111101100101", -- 8036 FREE #<CONS 0 8037>
 "00000000000000000001111101100110", -- 8037 FREE #<CONS 0 8038>
 "00000000000000000001111101100111", -- 8038 FREE #<CONS 0 8039>
 "00000000000000000001111101101000", -- 8039 FREE #<CONS 0 8040>
 "00000000000000000001111101101001", -- 8040 FREE #<CONS 0 8041>
 "00000000000000000001111101101010", -- 8041 FREE #<CONS 0 8042>
 "00000000000000000001111101101011", -- 8042 FREE #<CONS 0 8043>
 "00000000000000000001111101101100", -- 8043 FREE #<CONS 0 8044>
 "00000000000000000001111101101101", -- 8044 FREE #<CONS 0 8045>
 "00000000000000000001111101101110", -- 8045 FREE #<CONS 0 8046>
 "00000000000000000001111101101111", -- 8046 FREE #<CONS 0 8047>
 "00000000000000000001111101110000", -- 8047 FREE #<CONS 0 8048>
 "00000000000000000001111101110001", -- 8048 FREE #<CONS 0 8049>
 "00000000000000000001111101110010", -- 8049 FREE #<CONS 0 8050>
 "00000000000000000001111101110011", -- 8050 FREE #<CONS 0 8051>
 "00000000000000000001111101110100", -- 8051 FREE #<CONS 0 8052>
 "00000000000000000001111101110101", -- 8052 FREE #<CONS 0 8053>
 "00000000000000000001111101110110", -- 8053 FREE #<CONS 0 8054>
 "00000000000000000001111101110111", -- 8054 FREE #<CONS 0 8055>
 "00000000000000000001111101111000", -- 8055 FREE #<CONS 0 8056>
 "00000000000000000001111101111001", -- 8056 FREE #<CONS 0 8057>
 "00000000000000000001111101111010", -- 8057 FREE #<CONS 0 8058>
 "00000000000000000001111101111011", -- 8058 FREE #<CONS 0 8059>
 "00000000000000000001111101111100", -- 8059 FREE #<CONS 0 8060>
 "00000000000000000001111101111101", -- 8060 FREE #<CONS 0 8061>
 "00000000000000000001111101111110", -- 8061 FREE #<CONS 0 8062>
 "00000000000000000001111101111111", -- 8062 FREE #<CONS 0 8063>
 "00000000000000000001111110000000", -- 8063 FREE #<CONS 0 8064>
 "00000000000000000001111110000001", -- 8064 FREE #<CONS 0 8065>
 "00000000000000000001111110000010", -- 8065 FREE #<CONS 0 8066>
 "00000000000000000001111110000011", -- 8066 FREE #<CONS 0 8067>
 "00000000000000000001111110000100", -- 8067 FREE #<CONS 0 8068>
 "00000000000000000001111110000101", -- 8068 FREE #<CONS 0 8069>
 "00000000000000000001111110000110", -- 8069 FREE #<CONS 0 8070>
 "00000000000000000001111110000111", -- 8070 FREE #<CONS 0 8071>
 "00000000000000000001111110001000", -- 8071 FREE #<CONS 0 8072>
 "00000000000000000001111110001001", -- 8072 FREE #<CONS 0 8073>
 "00000000000000000001111110001010", -- 8073 FREE #<CONS 0 8074>
 "00000000000000000001111110001011", -- 8074 FREE #<CONS 0 8075>
 "00000000000000000001111110001100", -- 8075 FREE #<CONS 0 8076>
 "00000000000000000001111110001101", -- 8076 FREE #<CONS 0 8077>
 "00000000000000000001111110001110", -- 8077 FREE #<CONS 0 8078>
 "00000000000000000001111110001111", -- 8078 FREE #<CONS 0 8079>
 "00000000000000000001111110010000", -- 8079 FREE #<CONS 0 8080>
 "00000000000000000001111110010001", -- 8080 FREE #<CONS 0 8081>
 "00000000000000000001111110010010", -- 8081 FREE #<CONS 0 8082>
 "00000000000000000001111110010011", -- 8082 FREE #<CONS 0 8083>
 "00000000000000000001111110010100", -- 8083 FREE #<CONS 0 8084>
 "00000000000000000001111110010101", -- 8084 FREE #<CONS 0 8085>
 "00000000000000000001111110010110", -- 8085 FREE #<CONS 0 8086>
 "00000000000000000001111110010111", -- 8086 FREE #<CONS 0 8087>
 "00000000000000000001111110011000", -- 8087 FREE #<CONS 0 8088>
 "00000000000000000001111110011001", -- 8088 FREE #<CONS 0 8089>
 "00000000000000000001111110011010", -- 8089 FREE #<CONS 0 8090>
 "00000000000000000001111110011011", -- 8090 FREE #<CONS 0 8091>
 "00000000000000000001111110011100", -- 8091 FREE #<CONS 0 8092>
 "00000000000000000001111110011101", -- 8092 FREE #<CONS 0 8093>
 "00000000000000000001111110011110", -- 8093 FREE #<CONS 0 8094>
 "00000000000000000001111110011111", -- 8094 FREE #<CONS 0 8095>
 "00000000000000000001111110100000", -- 8095 FREE #<CONS 0 8096>
 "00000000000000000001111110100001", -- 8096 FREE #<CONS 0 8097>
 "00000000000000000001111110100010", -- 8097 FREE #<CONS 0 8098>
 "00000000000000000001111110100011", -- 8098 FREE #<CONS 0 8099>
 "00000000000000000001111110100100", -- 8099 FREE #<CONS 0 8100>
 "00000000000000000001111110100101", -- 8100 FREE #<CONS 0 8101>
 "00000000000000000001111110100110", -- 8101 FREE #<CONS 0 8102>
 "00000000000000000001111110100111", -- 8102 FREE #<CONS 0 8103>
 "00000000000000000001111110101000", -- 8103 FREE #<CONS 0 8104>
 "00000000000000000001111110101001", -- 8104 FREE #<CONS 0 8105>
 "00000000000000000001111110101010", -- 8105 FREE #<CONS 0 8106>
 "00000000000000000001111110101011", -- 8106 FREE #<CONS 0 8107>
 "00000000000000000001111110101100", -- 8107 FREE #<CONS 0 8108>
 "00000000000000000001111110101101", -- 8108 FREE #<CONS 0 8109>
 "00000000000000000001111110101110", -- 8109 FREE #<CONS 0 8110>
 "00000000000000000001111110101111", -- 8110 FREE #<CONS 0 8111>
 "00000000000000000001111110110000", -- 8111 FREE #<CONS 0 8112>
 "00000000000000000001111110110001", -- 8112 FREE #<CONS 0 8113>
 "00000000000000000001111110110010", -- 8113 FREE #<CONS 0 8114>
 "00000000000000000001111110110011", -- 8114 FREE #<CONS 0 8115>
 "00000000000000000001111110110100", -- 8115 FREE #<CONS 0 8116>
 "00000000000000000001111110110101", -- 8116 FREE #<CONS 0 8117>
 "00000000000000000001111110110110", -- 8117 FREE #<CONS 0 8118>
 "00000000000000000001111110110111", -- 8118 FREE #<CONS 0 8119>
 "00000000000000000001111110111000", -- 8119 FREE #<CONS 0 8120>
 "00000000000000000001111110111001", -- 8120 FREE #<CONS 0 8121>
 "00000000000000000001111110111010", -- 8121 FREE #<CONS 0 8122>
 "00000000000000000001111110111011", -- 8122 FREE #<CONS 0 8123>
 "00000000000000000001111110111100", -- 8123 FREE #<CONS 0 8124>
 "00000000000000000001111110111101", -- 8124 FREE #<CONS 0 8125>
 "00000000000000000001111110111110", -- 8125 FREE #<CONS 0 8126>
 "00000000000000000001111110111111", -- 8126 FREE #<CONS 0 8127>
 "00000000000000000001111111000000", -- 8127 FREE #<CONS 0 8128>
 "00000000000000000001111111000001", -- 8128 FREE #<CONS 0 8129>
 "00000000000000000001111111000010", -- 8129 FREE #<CONS 0 8130>
 "00000000000000000001111111000011", -- 8130 FREE #<CONS 0 8131>
 "00000000000000000001111111000100", -- 8131 FREE #<CONS 0 8132>
 "00000000000000000001111111000101", -- 8132 FREE #<CONS 0 8133>
 "00000000000000000001111111000110", -- 8133 FREE #<CONS 0 8134>
 "00000000000000000001111111000111", -- 8134 FREE #<CONS 0 8135>
 "00000000000000000001111111001000", -- 8135 FREE #<CONS 0 8136>
 "00000000000000000001111111001001", -- 8136 FREE #<CONS 0 8137>
 "00000000000000000001111111001010", -- 8137 FREE #<CONS 0 8138>
 "00000000000000000001111111001011", -- 8138 FREE #<CONS 0 8139>
 "00000000000000000001111111001100", -- 8139 FREE #<CONS 0 8140>
 "00000000000000000001111111001101", -- 8140 FREE #<CONS 0 8141>
 "00000000000000000001111111001110", -- 8141 FREE #<CONS 0 8142>
 "00000000000000000001111111001111", -- 8142 FREE #<CONS 0 8143>
 "00000000000000000001111111010000", -- 8143 FREE #<CONS 0 8144>
 "00000000000000000001111111010001", -- 8144 FREE #<CONS 0 8145>
 "00000000000000000001111111010010", -- 8145 FREE #<CONS 0 8146>
 "00000000000000000001111111010011", -- 8146 FREE #<CONS 0 8147>
 "00000000000000000001111111010100", -- 8147 FREE #<CONS 0 8148>
 "00000000000000000001111111010101", -- 8148 FREE #<CONS 0 8149>
 "00000000000000000001111111010110", -- 8149 FREE #<CONS 0 8150>
 "00000000000000000001111111010111", -- 8150 FREE #<CONS 0 8151>
 "00000000000000000001111111011000", -- 8151 FREE #<CONS 0 8152>
 "00000000000000000001111111011001", -- 8152 FREE #<CONS 0 8153>
 "00000000000000000001111111011010", -- 8153 FREE #<CONS 0 8154>
 "00000000000000000001111111011011", -- 8154 FREE #<CONS 0 8155>
 "00000000000000000001111111011100", -- 8155 FREE #<CONS 0 8156>
 "00000000000000000001111111011101", -- 8156 FREE #<CONS 0 8157>
 "00000000000000000001111111011110", -- 8157 FREE #<CONS 0 8158>
 "00000000000000000001111111011111", -- 8158 FREE #<CONS 0 8159>
 "00000000000000000001111111100000", -- 8159 FREE #<CONS 0 8160>
 "00000000000000000001111111100001", -- 8160 FREE #<CONS 0 8161>
 "00000000000000000001111111100010", -- 8161 FREE #<CONS 0 8162>
 "00000000000000000001111111100011", -- 8162 FREE #<CONS 0 8163>
 "00000000000000000001111111100100", -- 8163 FREE #<CONS 0 8164>
 "00000000000000000001111111100101", -- 8164 FREE #<CONS 0 8165>
 "00000000000000000001111111100110", -- 8165 FREE #<CONS 0 8166>
 "00000000000000000001111111100111", -- 8166 FREE #<CONS 0 8167>
 "00000000000000000001111111101000", -- 8167 FREE #<CONS 0 8168>
 "00000000000000000001111111101001", -- 8168 FREE #<CONS 0 8169>
 "00000000000000000001111111101010", -- 8169 FREE #<CONS 0 8170>
 "00000000000000000001111111101011", -- 8170 FREE #<CONS 0 8171>
 "00000000000000000001111111101100", -- 8171 FREE #<CONS 0 8172>
 "00000000000000000001111111101101", -- 8172 FREE #<CONS 0 8173>
 "00000000000000000001111111101110", -- 8173 FREE #<CONS 0 8174>
 "00000000000000000001111111101111", -- 8174 FREE #<CONS 0 8175>
 "00000000000000000001111111110000", -- 8175 FREE #<CONS 0 8176>
 "00000000000000000001111111110001", -- 8176 FREE #<CONS 0 8177>
 "00000000000000000001111111110010", -- 8177 FREE #<CONS 0 8178>
 "00000000000000000001111111110011", -- 8178 FREE #<CONS 0 8179>
 "00000000000000000001111111110100", -- 8179 FREE #<CONS 0 8180>
 "00000000000000000001111111110101", -- 8180 FREE #<CONS 0 8181>
 "00000000000000000001111111110110", -- 8181 FREE #<CONS 0 8182>
 "00000000000000000001111111110111", -- 8182 FREE #<CONS 0 8183>
 "00000000000000000001111111111000", -- 8183 FREE #<CONS 0 8184>
 "00000000000000000001111111111001", -- 8184 FREE #<CONS 0 8185>
 "00000000000000000001111111111010", -- 8185 FREE #<CONS 0 8186>
 "00000000000000000001111111111011", -- 8186 FREE #<CONS 0 8187>
 "00000000000000000001111111111100", -- 8187 FREE #<CONS 0 8188>
 "00000000000000000001111111111101", -- 8188 FREE #<CONS 0 8189>
 "00000000000000000001111111111110", -- 8189 FREE #<CONS 0 8190>
 "00000000000000000001111111111111", -- 8190 FREE #<CONS 0 8191>
 "00000000000000000010000000000000", -- 8191 FREE #<CONS 0 8192>
 "00000000000000000010000000000001", -- 8192 FREE #<CONS 0 8193>
 "00000000000000000010000000000010", -- 8193 FREE #<CONS 0 8194>
 "00000000000000000010000000000011", -- 8194 FREE #<CONS 0 8195>
 "00000000000000000010000000000100", -- 8195 FREE #<CONS 0 8196>
 "00000000000000000010000000000101", -- 8196 FREE #<CONS 0 8197>
 "00000000000000000010000000000110", -- 8197 FREE #<CONS 0 8198>
 "00000000000000000010000000000111", -- 8198 FREE #<CONS 0 8199>
 "00000000000000000010000000001000", -- 8199 FREE #<CONS 0 8200>
 "00000000000000000010000000001001", -- 8200 FREE #<CONS 0 8201>
 "00000000000000000010000000001010", -- 8201 FREE #<CONS 0 8202>
 "00000000000000000010000000001011", -- 8202 FREE #<CONS 0 8203>
 "00000000000000000010000000001100", -- 8203 FREE #<CONS 0 8204>
 "00000000000000000010000000001101", -- 8204 FREE #<CONS 0 8205>
 "00000000000000000010000000001110", -- 8205 FREE #<CONS 0 8206>
 "00000000000000000010000000001111", -- 8206 FREE #<CONS 0 8207>
 "00000000000000000010000000010000", -- 8207 FREE #<CONS 0 8208>
 "00000000000000000010000000010001", -- 8208 FREE #<CONS 0 8209>
 "00000000000000000010000000010010", -- 8209 FREE #<CONS 0 8210>
 "00000000000000000010000000010011", -- 8210 FREE #<CONS 0 8211>
 "00000000000000000010000000010100", -- 8211 FREE #<CONS 0 8212>
 "00000000000000000010000000010101", -- 8212 FREE #<CONS 0 8213>
 "00000000000000000010000000010110", -- 8213 FREE #<CONS 0 8214>
 "00000000000000000010000000010111", -- 8214 FREE #<CONS 0 8215>
 "00000000000000000010000000011000", -- 8215 FREE #<CONS 0 8216>
 "00000000000000000010000000011001", -- 8216 FREE #<CONS 0 8217>
 "00000000000000000010000000011010", -- 8217 FREE #<CONS 0 8218>
 "00000000000000000010000000011011", -- 8218 FREE #<CONS 0 8219>
 "00000000000000000010000000011100", -- 8219 FREE #<CONS 0 8220>
 "00000000000000000010000000011101", -- 8220 FREE #<CONS 0 8221>
 "00000000000000000010000000011110", -- 8221 FREE #<CONS 0 8222>
 "00000000000000000010000000011111", -- 8222 FREE #<CONS 0 8223>
 "00000000000000000010000000100000", -- 8223 FREE #<CONS 0 8224>
 "00000000000000000010000000100001", -- 8224 FREE #<CONS 0 8225>
 "00000000000000000010000000100010", -- 8225 FREE #<CONS 0 8226>
 "00000000000000000010000000100011", -- 8226 FREE #<CONS 0 8227>
 "00000000000000000010000000100100", -- 8227 FREE #<CONS 0 8228>
 "00000000000000000010000000100101", -- 8228 FREE #<CONS 0 8229>
 "00000000000000000010000000100110", -- 8229 FREE #<CONS 0 8230>
 "00000000000000000010000000100111", -- 8230 FREE #<CONS 0 8231>
 "00000000000000000010000000101000", -- 8231 FREE #<CONS 0 8232>
 "00000000000000000010000000101001", -- 8232 FREE #<CONS 0 8233>
 "00000000000000000010000000101010", -- 8233 FREE #<CONS 0 8234>
 "00000000000000000010000000101011", -- 8234 FREE #<CONS 0 8235>
 "00000000000000000010000000101100", -- 8235 FREE #<CONS 0 8236>
 "00000000000000000010000000101101", -- 8236 FREE #<CONS 0 8237>
 "00000000000000000010000000101110", -- 8237 FREE #<CONS 0 8238>
 "00000000000000000010000000101111", -- 8238 FREE #<CONS 0 8239>
 "00000000000000000010000000110000", -- 8239 FREE #<CONS 0 8240>
 "00000000000000000010000000110001", -- 8240 FREE #<CONS 0 8241>
 "00000000000000000010000000110010", -- 8241 FREE #<CONS 0 8242>
 "00000000000000000010000000110011", -- 8242 FREE #<CONS 0 8243>
 "00000000000000000010000000110100", -- 8243 FREE #<CONS 0 8244>
 "00000000000000000010000000110101", -- 8244 FREE #<CONS 0 8245>
 "00000000000000000010000000110110", -- 8245 FREE #<CONS 0 8246>
 "00000000000000000010000000110111", -- 8246 FREE #<CONS 0 8247>
 "00000000000000000010000000111000", -- 8247 FREE #<CONS 0 8248>
 "00000000000000000010000000111001", -- 8248 FREE #<CONS 0 8249>
 "00000000000000000010000000111010", -- 8249 FREE #<CONS 0 8250>
 "00000000000000000010000000111011", -- 8250 FREE #<CONS 0 8251>
 "00000000000000000010000000111100", -- 8251 FREE #<CONS 0 8252>
 "00000000000000000010000000111101", -- 8252 FREE #<CONS 0 8253>
 "00000000000000000010000000111110", -- 8253 FREE #<CONS 0 8254>
 "00000000000000000010000000111111", -- 8254 FREE #<CONS 0 8255>
 "00000000000000000010000001000000", -- 8255 FREE #<CONS 0 8256>
 "00000000000000000010000001000001", -- 8256 FREE #<CONS 0 8257>
 "00000000000000000010000001000010", -- 8257 FREE #<CONS 0 8258>
 "00000000000000000010000001000011", -- 8258 FREE #<CONS 0 8259>
 "00000000000000000010000001000100", -- 8259 FREE #<CONS 0 8260>
 "00000000000000000010000001000101", -- 8260 FREE #<CONS 0 8261>
 "00000000000000000010000001000110", -- 8261 FREE #<CONS 0 8262>
 "00000000000000000010000001000111", -- 8262 FREE #<CONS 0 8263>
 "00000000000000000010000001001000", -- 8263 FREE #<CONS 0 8264>
 "00000000000000000010000001001001", -- 8264 FREE #<CONS 0 8265>
 "00000000000000000010000001001010", -- 8265 FREE #<CONS 0 8266>
 "00000000000000000010000001001011", -- 8266 FREE #<CONS 0 8267>
 "00000000000000000010000001001100", -- 8267 FREE #<CONS 0 8268>
 "00000000000000000010000001001101", -- 8268 FREE #<CONS 0 8269>
 "00000000000000000010000001001110", -- 8269 FREE #<CONS 0 8270>
 "00000000000000000010000001001111", -- 8270 FREE #<CONS 0 8271>
 "00000000000000000010000001010000", -- 8271 FREE #<CONS 0 8272>
 "00000000000000000010000001010001", -- 8272 FREE #<CONS 0 8273>
 "00000000000000000010000001010010", -- 8273 FREE #<CONS 0 8274>
 "00000000000000000010000001010011", -- 8274 FREE #<CONS 0 8275>
 "00000000000000000010000001010100", -- 8275 FREE #<CONS 0 8276>
 "00000000000000000010000001010101", -- 8276 FREE #<CONS 0 8277>
 "00000000000000000010000001010110", -- 8277 FREE #<CONS 0 8278>
 "00000000000000000010000001010111", -- 8278 FREE #<CONS 0 8279>
 "00000000000000000010000001011000", -- 8279 FREE #<CONS 0 8280>
 "00000000000000000010000001011001", -- 8280 FREE #<CONS 0 8281>
 "00000000000000000010000001011010", -- 8281 FREE #<CONS 0 8282>
 "00000000000000000010000001011011", -- 8282 FREE #<CONS 0 8283>
 "00000000000000000010000001011100", -- 8283 FREE #<CONS 0 8284>
 "00000000000000000010000001011101", -- 8284 FREE #<CONS 0 8285>
 "00000000000000000010000001011110", -- 8285 FREE #<CONS 0 8286>
 "00000000000000000010000001011111", -- 8286 FREE #<CONS 0 8287>
 "00000000000000000010000001100000", -- 8287 FREE #<CONS 0 8288>
 "00000000000000000010000001100001", -- 8288 FREE #<CONS 0 8289>
 "00000000000000000010000001100010", -- 8289 FREE #<CONS 0 8290>
 "00000000000000000010000001100011", -- 8290 FREE #<CONS 0 8291>
 "00000000000000000010000001100100", -- 8291 FREE #<CONS 0 8292>
 "00000000000000000010000001100101", -- 8292 FREE #<CONS 0 8293>
 "00000000000000000010000001100110", -- 8293 FREE #<CONS 0 8294>
 "00000000000000000010000001100111", -- 8294 FREE #<CONS 0 8295>
 "00000000000000000010000001101000", -- 8295 FREE #<CONS 0 8296>
 "00000000000000000010000001101001", -- 8296 FREE #<CONS 0 8297>
 "00000000000000000010000001101010", -- 8297 FREE #<CONS 0 8298>
 "00000000000000000010000001101011", -- 8298 FREE #<CONS 0 8299>
 "00000000000000000010000001101100", -- 8299 FREE #<CONS 0 8300>
 "00000000000000000010000001101101", -- 8300 FREE #<CONS 0 8301>
 "00000000000000000010000001101110", -- 8301 FREE #<CONS 0 8302>
 "00000000000000000010000001101111", -- 8302 FREE #<CONS 0 8303>
 "00000000000000000010000001110000", -- 8303 FREE #<CONS 0 8304>
 "00000000000000000010000001110001", -- 8304 FREE #<CONS 0 8305>
 "00000000000000000010000001110010", -- 8305 FREE #<CONS 0 8306>
 "00000000000000000010000001110011", -- 8306 FREE #<CONS 0 8307>
 "00000000000000000010000001110100", -- 8307 FREE #<CONS 0 8308>
 "00000000000000000010000001110101", -- 8308 FREE #<CONS 0 8309>
 "00000000000000000010000001110110", -- 8309 FREE #<CONS 0 8310>
 "00000000000000000010000001110111", -- 8310 FREE #<CONS 0 8311>
 "00000000000000000010000001111000", -- 8311 FREE #<CONS 0 8312>
 "00000000000000000010000001111001", -- 8312 FREE #<CONS 0 8313>
 "00000000000000000010000001111010", -- 8313 FREE #<CONS 0 8314>
 "00000000000000000010000001111011", -- 8314 FREE #<CONS 0 8315>
 "00000000000000000010000001111100", -- 8315 FREE #<CONS 0 8316>
 "00000000000000000010000001111101", -- 8316 FREE #<CONS 0 8317>
 "00000000000000000010000001111110", -- 8317 FREE #<CONS 0 8318>
 "00000000000000000010000001111111", -- 8318 FREE #<CONS 0 8319>
 "00000000000000000010000010000000", -- 8319 FREE #<CONS 0 8320>
 "00000000000000000010000010000001", -- 8320 FREE #<CONS 0 8321>
 "00000000000000000010000010000010", -- 8321 FREE #<CONS 0 8322>
 "00000000000000000010000010000011", -- 8322 FREE #<CONS 0 8323>
 "00000000000000000010000010000100", -- 8323 FREE #<CONS 0 8324>
 "00000000000000000010000010000101", -- 8324 FREE #<CONS 0 8325>
 "00000000000000000010000010000110", -- 8325 FREE #<CONS 0 8326>
 "00000000000000000010000010000111", -- 8326 FREE #<CONS 0 8327>
 "00000000000000000010000010001000", -- 8327 FREE #<CONS 0 8328>
 "00000000000000000010000010001001", -- 8328 FREE #<CONS 0 8329>
 "00000000000000000010000010001010", -- 8329 FREE #<CONS 0 8330>
 "00000000000000000010000010001011", -- 8330 FREE #<CONS 0 8331>
 "00000000000000000010000010001100", -- 8331 FREE #<CONS 0 8332>
 "00000000000000000010000010001101", -- 8332 FREE #<CONS 0 8333>
 "00000000000000000010000010001110", -- 8333 FREE #<CONS 0 8334>
 "00000000000000000010000010001111", -- 8334 FREE #<CONS 0 8335>
 "00000000000000000010000010010000", -- 8335 FREE #<CONS 0 8336>
 "00000000000000000010000010010001", -- 8336 FREE #<CONS 0 8337>
 "00000000000000000010000010010010", -- 8337 FREE #<CONS 0 8338>
 "00000000000000000010000010010011", -- 8338 FREE #<CONS 0 8339>
 "00000000000000000010000010010100", -- 8339 FREE #<CONS 0 8340>
 "00000000000000000010000010010101", -- 8340 FREE #<CONS 0 8341>
 "00000000000000000010000010010110", -- 8341 FREE #<CONS 0 8342>
 "00000000000000000010000010010111", -- 8342 FREE #<CONS 0 8343>
 "00000000000000000010000010011000", -- 8343 FREE #<CONS 0 8344>
 "00000000000000000010000010011001", -- 8344 FREE #<CONS 0 8345>
 "00000000000000000010000010011010", -- 8345 FREE #<CONS 0 8346>
 "00000000000000000010000010011011", -- 8346 FREE #<CONS 0 8347>
 "00000000000000000010000010011100", -- 8347 FREE #<CONS 0 8348>
 "00000000000000000010000010011101", -- 8348 FREE #<CONS 0 8349>
 "00000000000000000010000010011110", -- 8349 FREE #<CONS 0 8350>
 "00000000000000000010000010011111", -- 8350 FREE #<CONS 0 8351>
 "00000000000000000010000010100000", -- 8351 FREE #<CONS 0 8352>
 "00000000000000000010000010100001", -- 8352 FREE #<CONS 0 8353>
 "00000000000000000010000010100010", -- 8353 FREE #<CONS 0 8354>
 "00000000000000000010000010100011", -- 8354 FREE #<CONS 0 8355>
 "00000000000000000010000010100100", -- 8355 FREE #<CONS 0 8356>
 "00000000000000000010000010100101", -- 8356 FREE #<CONS 0 8357>
 "00000000000000000010000010100110", -- 8357 FREE #<CONS 0 8358>
 "00000000000000000010000010100111", -- 8358 FREE #<CONS 0 8359>
 "00000000000000000010000010101000", -- 8359 FREE #<CONS 0 8360>
 "00000000000000000010000010101001", -- 8360 FREE #<CONS 0 8361>
 "00000000000000000010000010101010", -- 8361 FREE #<CONS 0 8362>
 "00000000000000000010000010101011", -- 8362 FREE #<CONS 0 8363>
 "00000000000000000010000010101100", -- 8363 FREE #<CONS 0 8364>
 "00000000000000000010000010101101", -- 8364 FREE #<CONS 0 8365>
 "00000000000000000010000010101110", -- 8365 FREE #<CONS 0 8366>
 "00000000000000000010000010101111", -- 8366 FREE #<CONS 0 8367>
 "00000000000000000010000010110000", -- 8367 FREE #<CONS 0 8368>
 "00000000000000000010000010110001", -- 8368 FREE #<CONS 0 8369>
 "00000000000000000010000010110010", -- 8369 FREE #<CONS 0 8370>
 "00000000000000000010000010110011", -- 8370 FREE #<CONS 0 8371>
 "00000000000000000010000010110100", -- 8371 FREE #<CONS 0 8372>
 "00000000000000000010000010110101", -- 8372 FREE #<CONS 0 8373>
 "00000000000000000010000010110110", -- 8373 FREE #<CONS 0 8374>
 "00000000000000000010000010110111", -- 8374 FREE #<CONS 0 8375>
 "00000000000000000010000010111000", -- 8375 FREE #<CONS 0 8376>
 "00000000000000000010000010111001", -- 8376 FREE #<CONS 0 8377>
 "00000000000000000010000010111010", -- 8377 FREE #<CONS 0 8378>
 "00000000000000000010000010111011", -- 8378 FREE #<CONS 0 8379>
 "00000000000000000010000010111100", -- 8379 FREE #<CONS 0 8380>
 "00000000000000000010000010111101", -- 8380 FREE #<CONS 0 8381>
 "00000000000000000010000010111110", -- 8381 FREE #<CONS 0 8382>
 "00000000000000000010000010111111", -- 8382 FREE #<CONS 0 8383>
 "00000000000000000010000011000000", -- 8383 FREE #<CONS 0 8384>
 "00000000000000000010000011000001", -- 8384 FREE #<CONS 0 8385>
 "00000000000000000010000011000010", -- 8385 FREE #<CONS 0 8386>
 "00000000000000000010000011000011", -- 8386 FREE #<CONS 0 8387>
 "00000000000000000010000011000100", -- 8387 FREE #<CONS 0 8388>
 "00000000000000000010000011000101", -- 8388 FREE #<CONS 0 8389>
 "00000000000000000010000011000110", -- 8389 FREE #<CONS 0 8390>
 "00000000000000000010000011000111", -- 8390 FREE #<CONS 0 8391>
 "00000000000000000010000011001000", -- 8391 FREE #<CONS 0 8392>
 "00000000000000000010000011001001", -- 8392 FREE #<CONS 0 8393>
 "00000000000000000010000011001010", -- 8393 FREE #<CONS 0 8394>
 "00000000000000000010000011001011", -- 8394 FREE #<CONS 0 8395>
 "00000000000000000010000011001100", -- 8395 FREE #<CONS 0 8396>
 "00000000000000000010000011001101", -- 8396 FREE #<CONS 0 8397>
 "00000000000000000010000011001110", -- 8397 FREE #<CONS 0 8398>
 "00000000000000000010000011001111", -- 8398 FREE #<CONS 0 8399>
 "00000000000000000010000011010000", -- 8399 FREE #<CONS 0 8400>
 "00000000000000000010000011010001", -- 8400 FREE #<CONS 0 8401>
 "00000000000000000010000011010010", -- 8401 FREE #<CONS 0 8402>
 "00000000000000000010000011010011", -- 8402 FREE #<CONS 0 8403>
 "00000000000000000010000011010100", -- 8403 FREE #<CONS 0 8404>
 "00000000000000000010000011010101", -- 8404 FREE #<CONS 0 8405>
 "00000000000000000010000011010110", -- 8405 FREE #<CONS 0 8406>
 "00000000000000000010000011010111", -- 8406 FREE #<CONS 0 8407>
 "00000000000000000010000011011000", -- 8407 FREE #<CONS 0 8408>
 "00000000000000000010000011011001", -- 8408 FREE #<CONS 0 8409>
 "00000000000000000010000011011010", -- 8409 FREE #<CONS 0 8410>
 "00000000000000000010000011011011", -- 8410 FREE #<CONS 0 8411>
 "00000000000000000010000011011100", -- 8411 FREE #<CONS 0 8412>
 "00000000000000000010000011011101", -- 8412 FREE #<CONS 0 8413>
 "00000000000000000010000011011110", -- 8413 FREE #<CONS 0 8414>
 "00000000000000000010000011011111", -- 8414 FREE #<CONS 0 8415>
 "00000000000000000010000011100000", -- 8415 FREE #<CONS 0 8416>
 "00000000000000000010000011100001", -- 8416 FREE #<CONS 0 8417>
 "00000000000000000010000011100010", -- 8417 FREE #<CONS 0 8418>
 "00000000000000000010000011100011", -- 8418 FREE #<CONS 0 8419>
 "00000000000000000010000011100100", -- 8419 FREE #<CONS 0 8420>
 "00000000000000000010000011100101", -- 8420 FREE #<CONS 0 8421>
 "00000000000000000010000011100110", -- 8421 FREE #<CONS 0 8422>
 "00000000000000000010000011100111", -- 8422 FREE #<CONS 0 8423>
 "00000000000000000010000011101000", -- 8423 FREE #<CONS 0 8424>
 "00000000000000000010000011101001", -- 8424 FREE #<CONS 0 8425>
 "00000000000000000010000011101010", -- 8425 FREE #<CONS 0 8426>
 "00000000000000000010000011101011", -- 8426 FREE #<CONS 0 8427>
 "00000000000000000010000011101100", -- 8427 FREE #<CONS 0 8428>
 "00000000000000000010000011101101", -- 8428 FREE #<CONS 0 8429>
 "00000000000000000010000011101110", -- 8429 FREE #<CONS 0 8430>
 "00000000000000000010000011101111", -- 8430 FREE #<CONS 0 8431>
 "00000000000000000010000011110000", -- 8431 FREE #<CONS 0 8432>
 "00000000000000000010000011110001", -- 8432 FREE #<CONS 0 8433>
 "00000000000000000010000011110010", -- 8433 FREE #<CONS 0 8434>
 "00000000000000000010000011110011", -- 8434 FREE #<CONS 0 8435>
 "00000000000000000010000011110100", -- 8435 FREE #<CONS 0 8436>
 "00000000000000000010000011110101", -- 8436 FREE #<CONS 0 8437>
 "00000000000000000010000011110110", -- 8437 FREE #<CONS 0 8438>
 "00000000000000000010000011110111", -- 8438 FREE #<CONS 0 8439>
 "00000000000000000010000011111000", -- 8439 FREE #<CONS 0 8440>
 "00000000000000000010000011111001", -- 8440 FREE #<CONS 0 8441>
 "00000000000000000010000011111010", -- 8441 FREE #<CONS 0 8442>
 "00000000000000000010000011111011", -- 8442 FREE #<CONS 0 8443>
 "00000000000000000010000011111100", -- 8443 FREE #<CONS 0 8444>
 "00000000000000000010000011111101", -- 8444 FREE #<CONS 0 8445>
 "00000000000000000010000011111110", -- 8445 FREE #<CONS 0 8446>
 "00000000000000000010000011111111", -- 8446 FREE #<CONS 0 8447>
 "00000000000000000010000100000000", -- 8447 FREE #<CONS 0 8448>
 "00000000000000000010000100000001", -- 8448 FREE #<CONS 0 8449>
 "00000000000000000010000100000010", -- 8449 FREE #<CONS 0 8450>
 "00000000000000000010000100000011", -- 8450 FREE #<CONS 0 8451>
 "00000000000000000010000100000100", -- 8451 FREE #<CONS 0 8452>
 "00000000000000000010000100000101", -- 8452 FREE #<CONS 0 8453>
 "00000000000000000010000100000110", -- 8453 FREE #<CONS 0 8454>
 "00000000000000000010000100000111", -- 8454 FREE #<CONS 0 8455>
 "00000000000000000010000100001000", -- 8455 FREE #<CONS 0 8456>
 "00000000000000000010000100001001", -- 8456 FREE #<CONS 0 8457>
 "00000000000000000010000100001010", -- 8457 FREE #<CONS 0 8458>
 "00000000000000000010000100001011", -- 8458 FREE #<CONS 0 8459>
 "00000000000000000010000100001100", -- 8459 FREE #<CONS 0 8460>
 "00000000000000000010000100001101", -- 8460 FREE #<CONS 0 8461>
 "00000000000000000010000100001110", -- 8461 FREE #<CONS 0 8462>
 "00000000000000000010000100001111", -- 8462 FREE #<CONS 0 8463>
 "00000000000000000010000100010000", -- 8463 FREE #<CONS 0 8464>
 "00000000000000000010000100010001", -- 8464 FREE #<CONS 0 8465>
 "00000000000000000010000100010010", -- 8465 FREE #<CONS 0 8466>
 "00000000000000000010000100010011", -- 8466 FREE #<CONS 0 8467>
 "00000000000000000010000100010100", -- 8467 FREE #<CONS 0 8468>
 "00000000000000000010000100010101", -- 8468 FREE #<CONS 0 8469>
 "00000000000000000010000100010110", -- 8469 FREE #<CONS 0 8470>
 "00000000000000000010000100010111", -- 8470 FREE #<CONS 0 8471>
 "00000000000000000010000100011000", -- 8471 FREE #<CONS 0 8472>
 "00000000000000000010000100011001", -- 8472 FREE #<CONS 0 8473>
 "00000000000000000010000100011010", -- 8473 FREE #<CONS 0 8474>
 "00000000000000000010000100011011", -- 8474 FREE #<CONS 0 8475>
 "00000000000000000010000100011100", -- 8475 FREE #<CONS 0 8476>
 "00000000000000000010000100011101", -- 8476 FREE #<CONS 0 8477>
 "00000000000000000010000100011110", -- 8477 FREE #<CONS 0 8478>
 "00000000000000000010000100011111", -- 8478 FREE #<CONS 0 8479>
 "00000000000000000010000100100000", -- 8479 FREE #<CONS 0 8480>
 "00000000000000000010000100100001", -- 8480 FREE #<CONS 0 8481>
 "00000000000000000010000100100010", -- 8481 FREE #<CONS 0 8482>
 "00000000000000000010000100100011", -- 8482 FREE #<CONS 0 8483>
 "00000000000000000010000100100100", -- 8483 FREE #<CONS 0 8484>
 "00000000000000000010000100100101", -- 8484 FREE #<CONS 0 8485>
 "00000000000000000010000100100110", -- 8485 FREE #<CONS 0 8486>
 "00000000000000000010000100100111", -- 8486 FREE #<CONS 0 8487>
 "00000000000000000010000100101000", -- 8487 FREE #<CONS 0 8488>
 "00000000000000000010000100101001", -- 8488 FREE #<CONS 0 8489>
 "00000000000000000010000100101010", -- 8489 FREE #<CONS 0 8490>
 "00000000000000000010000100101011", -- 8490 FREE #<CONS 0 8491>
 "00000000000000000010000100101100", -- 8491 FREE #<CONS 0 8492>
 "00000000000000000010000100101101", -- 8492 FREE #<CONS 0 8493>
 "00000000000000000010000100101110", -- 8493 FREE #<CONS 0 8494>
 "00000000000000000010000100101111", -- 8494 FREE #<CONS 0 8495>
 "00000000000000000010000100110000", -- 8495 FREE #<CONS 0 8496>
 "00000000000000000010000100110001", -- 8496 FREE #<CONS 0 8497>
 "00000000000000000010000100110010", -- 8497 FREE #<CONS 0 8498>
 "00000000000000000010000100110011", -- 8498 FREE #<CONS 0 8499>
 "00000000000000000010000100110100", -- 8499 FREE #<CONS 0 8500>
 "00000000000000000010000100110101", -- 8500 FREE #<CONS 0 8501>
 "00000000000000000010000100110110", -- 8501 FREE #<CONS 0 8502>
 "00000000000000000010000100110111", -- 8502 FREE #<CONS 0 8503>
 "00000000000000000010000100111000", -- 8503 FREE #<CONS 0 8504>
 "00000000000000000010000100111001", -- 8504 FREE #<CONS 0 8505>
 "00000000000000000010000100111010", -- 8505 FREE #<CONS 0 8506>
 "00000000000000000010000100111011", -- 8506 FREE #<CONS 0 8507>
 "00000000000000000010000100111100", -- 8507 FREE #<CONS 0 8508>
 "00000000000000000010000100111101", -- 8508 FREE #<CONS 0 8509>
 "00000000000000000010000100111110", -- 8509 FREE #<CONS 0 8510>
 "00000000000000000010000100111111", -- 8510 FREE #<CONS 0 8511>
 "00000000000000000010000101000000", -- 8511 FREE #<CONS 0 8512>
 "00000000000000000010000101000001", -- 8512 FREE #<CONS 0 8513>
 "00000000000000000010000101000010", -- 8513 FREE #<CONS 0 8514>
 "00000000000000000010000101000011", -- 8514 FREE #<CONS 0 8515>
 "00000000000000000010000101000100", -- 8515 FREE #<CONS 0 8516>
 "00000000000000000010000101000101", -- 8516 FREE #<CONS 0 8517>
 "00000000000000000010000101000110", -- 8517 FREE #<CONS 0 8518>
 "00000000000000000010000101000111", -- 8518 FREE #<CONS 0 8519>
 "00000000000000000010000101001000", -- 8519 FREE #<CONS 0 8520>
 "00000000000000000010000101001001", -- 8520 FREE #<CONS 0 8521>
 "00000000000000000010000101001010", -- 8521 FREE #<CONS 0 8522>
 "00000000000000000010000101001011", -- 8522 FREE #<CONS 0 8523>
 "00000000000000000010000101001100", -- 8523 FREE #<CONS 0 8524>
 "00000000000000000010000101001101", -- 8524 FREE #<CONS 0 8525>
 "00000000000000000010000101001110", -- 8525 FREE #<CONS 0 8526>
 "00000000000000000010000101001111", -- 8526 FREE #<CONS 0 8527>
 "00000000000000000010000101010000", -- 8527 FREE #<CONS 0 8528>
 "00000000000000000010000101010001", -- 8528 FREE #<CONS 0 8529>
 "00000000000000000010000101010010", -- 8529 FREE #<CONS 0 8530>
 "00000000000000000010000101010011", -- 8530 FREE #<CONS 0 8531>
 "00000000000000000010000101010100", -- 8531 FREE #<CONS 0 8532>
 "00000000000000000010000101010101", -- 8532 FREE #<CONS 0 8533>
 "00000000000000000010000101010110", -- 8533 FREE #<CONS 0 8534>
 "00000000000000000010000101010111", -- 8534 FREE #<CONS 0 8535>
 "00000000000000000010000101011000", -- 8535 FREE #<CONS 0 8536>
 "00000000000000000010000101011001", -- 8536 FREE #<CONS 0 8537>
 "00000000000000000010000101011010", -- 8537 FREE #<CONS 0 8538>
 "00000000000000000010000101011011", -- 8538 FREE #<CONS 0 8539>
 "00000000000000000010000101011100", -- 8539 FREE #<CONS 0 8540>
 "00000000000000000010000101011101", -- 8540 FREE #<CONS 0 8541>
 "00000000000000000010000101011110", -- 8541 FREE #<CONS 0 8542>
 "00000000000000000010000101011111", -- 8542 FREE #<CONS 0 8543>
 "00000000000000000010000101100000", -- 8543 FREE #<CONS 0 8544>
 "00000000000000000010000101100001", -- 8544 FREE #<CONS 0 8545>
 "00000000000000000010000101100010", -- 8545 FREE #<CONS 0 8546>
 "00000000000000000010000101100011", -- 8546 FREE #<CONS 0 8547>
 "00000000000000000010000101100100", -- 8547 FREE #<CONS 0 8548>
 "00000000000000000010000101100101", -- 8548 FREE #<CONS 0 8549>
 "00000000000000000010000101100110", -- 8549 FREE #<CONS 0 8550>
 "00000000000000000010000101100111", -- 8550 FREE #<CONS 0 8551>
 "00000000000000000010000101101000", -- 8551 FREE #<CONS 0 8552>
 "00000000000000000010000101101001", -- 8552 FREE #<CONS 0 8553>
 "00000000000000000010000101101010", -- 8553 FREE #<CONS 0 8554>
 "00000000000000000010000101101011", -- 8554 FREE #<CONS 0 8555>
 "00000000000000000010000101101100", -- 8555 FREE #<CONS 0 8556>
 "00000000000000000010000101101101", -- 8556 FREE #<CONS 0 8557>
 "00000000000000000010000101101110", -- 8557 FREE #<CONS 0 8558>
 "00000000000000000010000101101111", -- 8558 FREE #<CONS 0 8559>
 "00000000000000000010000101110000", -- 8559 FREE #<CONS 0 8560>
 "00000000000000000010000101110001", -- 8560 FREE #<CONS 0 8561>
 "00000000000000000010000101110010", -- 8561 FREE #<CONS 0 8562>
 "00000000000000000010000101110011", -- 8562 FREE #<CONS 0 8563>
 "00000000000000000010000101110100", -- 8563 FREE #<CONS 0 8564>
 "00000000000000000010000101110101", -- 8564 FREE #<CONS 0 8565>
 "00000000000000000010000101110110", -- 8565 FREE #<CONS 0 8566>
 "00000000000000000010000101110111", -- 8566 FREE #<CONS 0 8567>
 "00000000000000000010000101111000", -- 8567 FREE #<CONS 0 8568>
 "00000000000000000010000101111001", -- 8568 FREE #<CONS 0 8569>
 "00000000000000000010000101111010", -- 8569 FREE #<CONS 0 8570>
 "00000000000000000010000101111011", -- 8570 FREE #<CONS 0 8571>
 "00000000000000000010000101111100", -- 8571 FREE #<CONS 0 8572>
 "00000000000000000010000101111101", -- 8572 FREE #<CONS 0 8573>
 "00000000000000000010000101111110", -- 8573 FREE #<CONS 0 8574>
 "00000000000000000010000101111111", -- 8574 FREE #<CONS 0 8575>
 "00000000000000000010000110000000", -- 8575 FREE #<CONS 0 8576>
 "00000000000000000010000110000001", -- 8576 FREE #<CONS 0 8577>
 "00000000000000000010000110000010", -- 8577 FREE #<CONS 0 8578>
 "00000000000000000010000110000011", -- 8578 FREE #<CONS 0 8579>
 "00000000000000000010000110000100", -- 8579 FREE #<CONS 0 8580>
 "00000000000000000010000110000101", -- 8580 FREE #<CONS 0 8581>
 "00000000000000000010000110000110", -- 8581 FREE #<CONS 0 8582>
 "00000000000000000010000110000111", -- 8582 FREE #<CONS 0 8583>
 "00000000000000000010000110001000", -- 8583 FREE #<CONS 0 8584>
 "00000000000000000010000110001001", -- 8584 FREE #<CONS 0 8585>
 "00000000000000000010000110001010", -- 8585 FREE #<CONS 0 8586>
 "00000000000000000010000110001011", -- 8586 FREE #<CONS 0 8587>
 "00000000000000000010000110001100", -- 8587 FREE #<CONS 0 8588>
 "00000000000000000010000110001101", -- 8588 FREE #<CONS 0 8589>
 "00000000000000000010000110001110", -- 8589 FREE #<CONS 0 8590>
 "00000000000000000010000110001111", -- 8590 FREE #<CONS 0 8591>
 "00000000000000000010000110010000", -- 8591 FREE #<CONS 0 8592>
 "00000000000000000010000110010001", -- 8592 FREE #<CONS 0 8593>
 "00000000000000000010000110010010", -- 8593 FREE #<CONS 0 8594>
 "00000000000000000010000110010011", -- 8594 FREE #<CONS 0 8595>
 "00000000000000000010000110010100", -- 8595 FREE #<CONS 0 8596>
 "00000000000000000010000110010101", -- 8596 FREE #<CONS 0 8597>
 "00000000000000000010000110010110", -- 8597 FREE #<CONS 0 8598>
 "00000000000000000010000110010111", -- 8598 FREE #<CONS 0 8599>
 "00000000000000000010000110011000", -- 8599 FREE #<CONS 0 8600>
 "00000000000000000010000110011001", -- 8600 FREE #<CONS 0 8601>
 "00000000000000000010000110011010", -- 8601 FREE #<CONS 0 8602>
 "00000000000000000010000110011011", -- 8602 FREE #<CONS 0 8603>
 "00000000000000000010000110011100", -- 8603 FREE #<CONS 0 8604>
 "00000000000000000010000110011101", -- 8604 FREE #<CONS 0 8605>
 "00000000000000000010000110011110", -- 8605 FREE #<CONS 0 8606>
 "00000000000000000010000110011111", -- 8606 FREE #<CONS 0 8607>
 "00000000000000000010000110100000", -- 8607 FREE #<CONS 0 8608>
 "00000000000000000010000110100001", -- 8608 FREE #<CONS 0 8609>
 "00000000000000000010000110100010", -- 8609 FREE #<CONS 0 8610>
 "00000000000000000010000110100011", -- 8610 FREE #<CONS 0 8611>
 "00000000000000000010000110100100", -- 8611 FREE #<CONS 0 8612>
 "00000000000000000010000110100101", -- 8612 FREE #<CONS 0 8613>
 "00000000000000000010000110100110", -- 8613 FREE #<CONS 0 8614>
 "00000000000000000010000110100111", -- 8614 FREE #<CONS 0 8615>
 "00000000000000000010000110101000", -- 8615 FREE #<CONS 0 8616>
 "00000000000000000010000110101001", -- 8616 FREE #<CONS 0 8617>
 "00000000000000000010000110101010", -- 8617 FREE #<CONS 0 8618>
 "00000000000000000010000110101011", -- 8618 FREE #<CONS 0 8619>
 "00000000000000000010000110101100", -- 8619 FREE #<CONS 0 8620>
 "00000000000000000010000110101101", -- 8620 FREE #<CONS 0 8621>
 "00000000000000000010000110101110", -- 8621 FREE #<CONS 0 8622>
 "00000000000000000010000110101111", -- 8622 FREE #<CONS 0 8623>
 "00000000000000000010000110110000", -- 8623 FREE #<CONS 0 8624>
 "00000000000000000010000110110001", -- 8624 FREE #<CONS 0 8625>
 "00000000000000000010000110110010", -- 8625 FREE #<CONS 0 8626>
 "00000000000000000010000110110011", -- 8626 FREE #<CONS 0 8627>
 "00000000000000000010000110110100", -- 8627 FREE #<CONS 0 8628>
 "00000000000000000010000110110101", -- 8628 FREE #<CONS 0 8629>
 "00000000000000000010000110110110", -- 8629 FREE #<CONS 0 8630>
 "00000000000000000010000110110111", -- 8630 FREE #<CONS 0 8631>
 "00000000000000000010000110111000", -- 8631 FREE #<CONS 0 8632>
 "00000000000000000010000110111001", -- 8632 FREE #<CONS 0 8633>
 "00000000000000000010000110111010", -- 8633 FREE #<CONS 0 8634>
 "00000000000000000010000110111011", -- 8634 FREE #<CONS 0 8635>
 "00000000000000000010000110111100", -- 8635 FREE #<CONS 0 8636>
 "00000000000000000010000110111101", -- 8636 FREE #<CONS 0 8637>
 "00000000000000000010000110111110", -- 8637 FREE #<CONS 0 8638>
 "00000000000000000010000110111111", -- 8638 FREE #<CONS 0 8639>
 "00000000000000000010000111000000", -- 8639 FREE #<CONS 0 8640>
 "00000000000000000010000111000001", -- 8640 FREE #<CONS 0 8641>
 "00000000000000000010000111000010", -- 8641 FREE #<CONS 0 8642>
 "00000000000000000010000111000011", -- 8642 FREE #<CONS 0 8643>
 "00000000000000000010000111000100", -- 8643 FREE #<CONS 0 8644>
 "00000000000000000010000111000101", -- 8644 FREE #<CONS 0 8645>
 "00000000000000000010000111000110", -- 8645 FREE #<CONS 0 8646>
 "00000000000000000010000111000111", -- 8646 FREE #<CONS 0 8647>
 "00000000000000000010000111001000", -- 8647 FREE #<CONS 0 8648>
 "00000000000000000010000111001001", -- 8648 FREE #<CONS 0 8649>
 "00000000000000000010000111001010", -- 8649 FREE #<CONS 0 8650>
 "00000000000000000010000111001011", -- 8650 FREE #<CONS 0 8651>
 "00000000000000000010000111001100", -- 8651 FREE #<CONS 0 8652>
 "00000000000000000010000111001101", -- 8652 FREE #<CONS 0 8653>
 "00000000000000000010000111001110", -- 8653 FREE #<CONS 0 8654>
 "00000000000000000010000111001111", -- 8654 FREE #<CONS 0 8655>
 "00000000000000000010000111010000", -- 8655 FREE #<CONS 0 8656>
 "00000000000000000010000111010001", -- 8656 FREE #<CONS 0 8657>
 "00000000000000000010000111010010", -- 8657 FREE #<CONS 0 8658>
 "00000000000000000010000111010011", -- 8658 FREE #<CONS 0 8659>
 "00000000000000000010000111010100", -- 8659 FREE #<CONS 0 8660>
 "00000000000000000010000111010101", -- 8660 FREE #<CONS 0 8661>
 "00000000000000000010000111010110", -- 8661 FREE #<CONS 0 8662>
 "00000000000000000010000111010111", -- 8662 FREE #<CONS 0 8663>
 "00000000000000000010000111011000", -- 8663 FREE #<CONS 0 8664>
 "00000000000000000010000111011001", -- 8664 FREE #<CONS 0 8665>
 "00000000000000000010000111011010", -- 8665 FREE #<CONS 0 8666>
 "00000000000000000010000111011011", -- 8666 FREE #<CONS 0 8667>
 "00000000000000000010000111011100", -- 8667 FREE #<CONS 0 8668>
 "00000000000000000010000111011101", -- 8668 FREE #<CONS 0 8669>
 "00000000000000000010000111011110", -- 8669 FREE #<CONS 0 8670>
 "00000000000000000010000111011111", -- 8670 FREE #<CONS 0 8671>
 "00000000000000000010000111100000", -- 8671 FREE #<CONS 0 8672>
 "00000000000000000010000111100001", -- 8672 FREE #<CONS 0 8673>
 "00000000000000000010000111100010", -- 8673 FREE #<CONS 0 8674>
 "00000000000000000010000111100011", -- 8674 FREE #<CONS 0 8675>
 "00000000000000000010000111100100", -- 8675 FREE #<CONS 0 8676>
 "00000000000000000010000111100101", -- 8676 FREE #<CONS 0 8677>
 "00000000000000000010000111100110", -- 8677 FREE #<CONS 0 8678>
 "00000000000000000010000111100111", -- 8678 FREE #<CONS 0 8679>
 "00000000000000000010000111101000", -- 8679 FREE #<CONS 0 8680>
 "00000000000000000010000111101001", -- 8680 FREE #<CONS 0 8681>
 "00000000000000000010000111101010", -- 8681 FREE #<CONS 0 8682>
 "00000000000000000010000111101011", -- 8682 FREE #<CONS 0 8683>
 "00000000000000000010000111101100", -- 8683 FREE #<CONS 0 8684>
 "00000000000000000010000111101101", -- 8684 FREE #<CONS 0 8685>
 "00000000000000000010000111101110", -- 8685 FREE #<CONS 0 8686>
 "00000000000000000010000111101111", -- 8686 FREE #<CONS 0 8687>
 "00000000000000000010000111110000", -- 8687 FREE #<CONS 0 8688>
 "00000000000000000010000111110001", -- 8688 FREE #<CONS 0 8689>
 "00000000000000000010000111110010", -- 8689 FREE #<CONS 0 8690>
 "00000000000000000010000111110011", -- 8690 FREE #<CONS 0 8691>
 "00000000000000000010000111110100", -- 8691 FREE #<CONS 0 8692>
 "00000000000000000010000111110101", -- 8692 FREE #<CONS 0 8693>
 "00000000000000000010000111110110", -- 8693 FREE #<CONS 0 8694>
 "00000000000000000010000111110111", -- 8694 FREE #<CONS 0 8695>
 "00000000000000000010000111111000", -- 8695 FREE #<CONS 0 8696>
 "00000000000000000010000111111001", -- 8696 FREE #<CONS 0 8697>
 "00000000000000000010000111111010", -- 8697 FREE #<CONS 0 8698>
 "00000000000000000010000111111011", -- 8698 FREE #<CONS 0 8699>
 "00000000000000000010000111111100", -- 8699 FREE #<CONS 0 8700>
 "00000000000000000010000111111101", -- 8700 FREE #<CONS 0 8701>
 "00000000000000000010000111111110", -- 8701 FREE #<CONS 0 8702>
 "00000000000000000010000111111111", -- 8702 FREE #<CONS 0 8703>
 "00000000000000000010001000000000", -- 8703 FREE #<CONS 0 8704>
 "00000000000000000010001000000001", -- 8704 FREE #<CONS 0 8705>
 "00000000000000000010001000000010", -- 8705 FREE #<CONS 0 8706>
 "00000000000000000010001000000011", -- 8706 FREE #<CONS 0 8707>
 "00000000000000000010001000000100", -- 8707 FREE #<CONS 0 8708>
 "00000000000000000010001000000101", -- 8708 FREE #<CONS 0 8709>
 "00000000000000000010001000000110", -- 8709 FREE #<CONS 0 8710>
 "00000000000000000010001000000111", -- 8710 FREE #<CONS 0 8711>
 "00000000000000000010001000001000", -- 8711 FREE #<CONS 0 8712>
 "00000000000000000010001000001001", -- 8712 FREE #<CONS 0 8713>
 "00000000000000000010001000001010", -- 8713 FREE #<CONS 0 8714>
 "00000000000000000010001000001011", -- 8714 FREE #<CONS 0 8715>
 "00000000000000000010001000001100", -- 8715 FREE #<CONS 0 8716>
 "00000000000000000010001000001101", -- 8716 FREE #<CONS 0 8717>
 "00000000000000000010001000001110", -- 8717 FREE #<CONS 0 8718>
 "00000000000000000010001000001111", -- 8718 FREE #<CONS 0 8719>
 "00000000000000000010001000010000", -- 8719 FREE #<CONS 0 8720>
 "00000000000000000010001000010001", -- 8720 FREE #<CONS 0 8721>
 "00000000000000000010001000010010", -- 8721 FREE #<CONS 0 8722>
 "00000000000000000010001000010011", -- 8722 FREE #<CONS 0 8723>
 "00000000000000000010001000010100", -- 8723 FREE #<CONS 0 8724>
 "00000000000000000010001000010101", -- 8724 FREE #<CONS 0 8725>
 "00000000000000000010001000010110", -- 8725 FREE #<CONS 0 8726>
 "00000000000000000010001000010111", -- 8726 FREE #<CONS 0 8727>
 "00000000000000000010001000011000", -- 8727 FREE #<CONS 0 8728>
 "00000000000000000010001000011001", -- 8728 FREE #<CONS 0 8729>
 "00000000000000000010001000011010", -- 8729 FREE #<CONS 0 8730>
 "00000000000000000010001000011011", -- 8730 FREE #<CONS 0 8731>
 "00000000000000000010001000011100", -- 8731 FREE #<CONS 0 8732>
 "00000000000000000010001000011101", -- 8732 FREE #<CONS 0 8733>
 "00000000000000000010001000011110", -- 8733 FREE #<CONS 0 8734>
 "00000000000000000010001000011111", -- 8734 FREE #<CONS 0 8735>
 "00000000000000000010001000100000", -- 8735 FREE #<CONS 0 8736>
 "00000000000000000010001000100001", -- 8736 FREE #<CONS 0 8737>
 "00000000000000000010001000100010", -- 8737 FREE #<CONS 0 8738>
 "00000000000000000010001000100011", -- 8738 FREE #<CONS 0 8739>
 "00000000000000000010001000100100", -- 8739 FREE #<CONS 0 8740>
 "00000000000000000010001000100101", -- 8740 FREE #<CONS 0 8741>
 "00000000000000000010001000100110", -- 8741 FREE #<CONS 0 8742>
 "00000000000000000010001000100111", -- 8742 FREE #<CONS 0 8743>
 "00000000000000000010001000101000", -- 8743 FREE #<CONS 0 8744>
 "00000000000000000010001000101001", -- 8744 FREE #<CONS 0 8745>
 "00000000000000000010001000101010", -- 8745 FREE #<CONS 0 8746>
 "00000000000000000010001000101011", -- 8746 FREE #<CONS 0 8747>
 "00000000000000000010001000101100", -- 8747 FREE #<CONS 0 8748>
 "00000000000000000010001000101101", -- 8748 FREE #<CONS 0 8749>
 "00000000000000000010001000101110", -- 8749 FREE #<CONS 0 8750>
 "00000000000000000010001000101111", -- 8750 FREE #<CONS 0 8751>
 "00000000000000000010001000110000", -- 8751 FREE #<CONS 0 8752>
 "00000000000000000010001000110001", -- 8752 FREE #<CONS 0 8753>
 "00000000000000000010001000110010", -- 8753 FREE #<CONS 0 8754>
 "00000000000000000010001000110011", -- 8754 FREE #<CONS 0 8755>
 "00000000000000000010001000110100", -- 8755 FREE #<CONS 0 8756>
 "00000000000000000010001000110101", -- 8756 FREE #<CONS 0 8757>
 "00000000000000000010001000110110", -- 8757 FREE #<CONS 0 8758>
 "00000000000000000010001000110111", -- 8758 FREE #<CONS 0 8759>
 "00000000000000000010001000111000", -- 8759 FREE #<CONS 0 8760>
 "00000000000000000010001000111001", -- 8760 FREE #<CONS 0 8761>
 "00000000000000000010001000111010", -- 8761 FREE #<CONS 0 8762>
 "00000000000000000010001000111011", -- 8762 FREE #<CONS 0 8763>
 "00000000000000000010001000111100", -- 8763 FREE #<CONS 0 8764>
 "00000000000000000010001000111101", -- 8764 FREE #<CONS 0 8765>
 "00000000000000000010001000111110", -- 8765 FREE #<CONS 0 8766>
 "00000000000000000010001000111111", -- 8766 FREE #<CONS 0 8767>
 "00000000000000000010001001000000", -- 8767 FREE #<CONS 0 8768>
 "00000000000000000010001001000001", -- 8768 FREE #<CONS 0 8769>
 "00000000000000000010001001000010", -- 8769 FREE #<CONS 0 8770>
 "00000000000000000010001001000011", -- 8770 FREE #<CONS 0 8771>
 "00000000000000000010001001000100", -- 8771 FREE #<CONS 0 8772>
 "00000000000000000010001001000101", -- 8772 FREE #<CONS 0 8773>
 "00000000000000000010001001000110", -- 8773 FREE #<CONS 0 8774>
 "00000000000000000010001001000111", -- 8774 FREE #<CONS 0 8775>
 "00000000000000000010001001001000", -- 8775 FREE #<CONS 0 8776>
 "00000000000000000010001001001001", -- 8776 FREE #<CONS 0 8777>
 "00000000000000000010001001001010", -- 8777 FREE #<CONS 0 8778>
 "00000000000000000010001001001011", -- 8778 FREE #<CONS 0 8779>
 "00000000000000000010001001001100", -- 8779 FREE #<CONS 0 8780>
 "00000000000000000010001001001101", -- 8780 FREE #<CONS 0 8781>
 "00000000000000000010001001001110", -- 8781 FREE #<CONS 0 8782>
 "00000000000000000010001001001111", -- 8782 FREE #<CONS 0 8783>
 "00000000000000000010001001010000", -- 8783 FREE #<CONS 0 8784>
 "00000000000000000010001001010001", -- 8784 FREE #<CONS 0 8785>
 "00000000000000000010001001010010", -- 8785 FREE #<CONS 0 8786>
 "00000000000000000010001001010011", -- 8786 FREE #<CONS 0 8787>
 "00000000000000000010001001010100", -- 8787 FREE #<CONS 0 8788>
 "00000000000000000010001001010101", -- 8788 FREE #<CONS 0 8789>
 "00000000000000000010001001010110", -- 8789 FREE #<CONS 0 8790>
 "00000000000000000010001001010111", -- 8790 FREE #<CONS 0 8791>
 "00000000000000000010001001011000", -- 8791 FREE #<CONS 0 8792>
 "00000000000000000010001001011001", -- 8792 FREE #<CONS 0 8793>
 "00000000000000000010001001011010", -- 8793 FREE #<CONS 0 8794>
 "00000000000000000010001001011011", -- 8794 FREE #<CONS 0 8795>
 "00000000000000000010001001011100", -- 8795 FREE #<CONS 0 8796>
 "00000000000000000010001001011101", -- 8796 FREE #<CONS 0 8797>
 "00000000000000000010001001011110", -- 8797 FREE #<CONS 0 8798>
 "00000000000000000010001001011111", -- 8798 FREE #<CONS 0 8799>
 "00000000000000000010001001100000", -- 8799 FREE #<CONS 0 8800>
 "00000000000000000010001001100001", -- 8800 FREE #<CONS 0 8801>
 "00000000000000000010001001100010", -- 8801 FREE #<CONS 0 8802>
 "00000000000000000010001001100011", -- 8802 FREE #<CONS 0 8803>
 "00000000000000000010001001100100", -- 8803 FREE #<CONS 0 8804>
 "00000000000000000010001001100101", -- 8804 FREE #<CONS 0 8805>
 "00000000000000000010001001100110", -- 8805 FREE #<CONS 0 8806>
 "00000000000000000010001001100111", -- 8806 FREE #<CONS 0 8807>
 "00000000000000000010001001101000", -- 8807 FREE #<CONS 0 8808>
 "00000000000000000010001001101001", -- 8808 FREE #<CONS 0 8809>
 "00000000000000000010001001101010", -- 8809 FREE #<CONS 0 8810>
 "00000000000000000010001001101011", -- 8810 FREE #<CONS 0 8811>
 "00000000000000000010001001101100", -- 8811 FREE #<CONS 0 8812>
 "00000000000000000010001001101101", -- 8812 FREE #<CONS 0 8813>
 "00000000000000000010001001101110", -- 8813 FREE #<CONS 0 8814>
 "00000000000000000010001001101111", -- 8814 FREE #<CONS 0 8815>
 "00000000000000000010001001110000", -- 8815 FREE #<CONS 0 8816>
 "00000000000000000010001001110001", -- 8816 FREE #<CONS 0 8817>
 "00000000000000000010001001110010", -- 8817 FREE #<CONS 0 8818>
 "00000000000000000010001001110011", -- 8818 FREE #<CONS 0 8819>
 "00000000000000000010001001110100", -- 8819 FREE #<CONS 0 8820>
 "00000000000000000010001001110101", -- 8820 FREE #<CONS 0 8821>
 "00000000000000000010001001110110", -- 8821 FREE #<CONS 0 8822>
 "00000000000000000010001001110111", -- 8822 FREE #<CONS 0 8823>
 "00000000000000000010001001111000", -- 8823 FREE #<CONS 0 8824>
 "00000000000000000010001001111001", -- 8824 FREE #<CONS 0 8825>
 "00000000000000000010001001111010", -- 8825 FREE #<CONS 0 8826>
 "00000000000000000010001001111011", -- 8826 FREE #<CONS 0 8827>
 "00000000000000000010001001111100", -- 8827 FREE #<CONS 0 8828>
 "00000000000000000010001001111101", -- 8828 FREE #<CONS 0 8829>
 "00000000000000000010001001111110", -- 8829 FREE #<CONS 0 8830>
 "00000000000000000010001001111111", -- 8830 FREE #<CONS 0 8831>
 "00000000000000000010001010000000", -- 8831 FREE #<CONS 0 8832>
 "00000000000000000010001010000001", -- 8832 FREE #<CONS 0 8833>
 "00000000000000000010001010000010", -- 8833 FREE #<CONS 0 8834>
 "00000000000000000010001010000011", -- 8834 FREE #<CONS 0 8835>
 "00000000000000000010001010000100", -- 8835 FREE #<CONS 0 8836>
 "00000000000000000010001010000101", -- 8836 FREE #<CONS 0 8837>
 "00000000000000000010001010000110", -- 8837 FREE #<CONS 0 8838>
 "00000000000000000010001010000111", -- 8838 FREE #<CONS 0 8839>
 "00000000000000000010001010001000", -- 8839 FREE #<CONS 0 8840>
 "00000000000000000010001010001001", -- 8840 FREE #<CONS 0 8841>
 "00000000000000000010001010001010", -- 8841 FREE #<CONS 0 8842>
 "00000000000000000010001010001011", -- 8842 FREE #<CONS 0 8843>
 "00000000000000000010001010001100", -- 8843 FREE #<CONS 0 8844>
 "00000000000000000010001010001101", -- 8844 FREE #<CONS 0 8845>
 "00000000000000000010001010001110", -- 8845 FREE #<CONS 0 8846>
 "00000000000000000010001010001111", -- 8846 FREE #<CONS 0 8847>
 "00000000000000000010001010010000", -- 8847 FREE #<CONS 0 8848>
 "00000000000000000010001010010001", -- 8848 FREE #<CONS 0 8849>
 "00000000000000000010001010010010", -- 8849 FREE #<CONS 0 8850>
 "00000000000000000010001010010011", -- 8850 FREE #<CONS 0 8851>
 "00000000000000000010001010010100", -- 8851 FREE #<CONS 0 8852>
 "00000000000000000010001010010101", -- 8852 FREE #<CONS 0 8853>
 "00000000000000000010001010010110", -- 8853 FREE #<CONS 0 8854>
 "00000000000000000010001010010111", -- 8854 FREE #<CONS 0 8855>
 "00000000000000000010001010011000", -- 8855 FREE #<CONS 0 8856>
 "00000000000000000010001010011001", -- 8856 FREE #<CONS 0 8857>
 "00000000000000000010001010011010", -- 8857 FREE #<CONS 0 8858>
 "00000000000000000010001010011011", -- 8858 FREE #<CONS 0 8859>
 "00000000000000000010001010011100", -- 8859 FREE #<CONS 0 8860>
 "00000000000000000010001010011101", -- 8860 FREE #<CONS 0 8861>
 "00000000000000000010001010011110", -- 8861 FREE #<CONS 0 8862>
 "00000000000000000010001010011111", -- 8862 FREE #<CONS 0 8863>
 "00000000000000000010001010100000", -- 8863 FREE #<CONS 0 8864>
 "00000000000000000010001010100001", -- 8864 FREE #<CONS 0 8865>
 "00000000000000000010001010100010", -- 8865 FREE #<CONS 0 8866>
 "00000000000000000010001010100011", -- 8866 FREE #<CONS 0 8867>
 "00000000000000000010001010100100", -- 8867 FREE #<CONS 0 8868>
 "00000000000000000010001010100101", -- 8868 FREE #<CONS 0 8869>
 "00000000000000000010001010100110", -- 8869 FREE #<CONS 0 8870>
 "00000000000000000010001010100111", -- 8870 FREE #<CONS 0 8871>
 "00000000000000000010001010101000", -- 8871 FREE #<CONS 0 8872>
 "00000000000000000010001010101001", -- 8872 FREE #<CONS 0 8873>
 "00000000000000000010001010101010", -- 8873 FREE #<CONS 0 8874>
 "00000000000000000010001010101011", -- 8874 FREE #<CONS 0 8875>
 "00000000000000000010001010101100", -- 8875 FREE #<CONS 0 8876>
 "00000000000000000010001010101101", -- 8876 FREE #<CONS 0 8877>
 "00000000000000000010001010101110", -- 8877 FREE #<CONS 0 8878>
 "00000000000000000010001010101111", -- 8878 FREE #<CONS 0 8879>
 "00000000000000000010001010110000", -- 8879 FREE #<CONS 0 8880>
 "00000000000000000010001010110001", -- 8880 FREE #<CONS 0 8881>
 "00000000000000000010001010110010", -- 8881 FREE #<CONS 0 8882>
 "00000000000000000010001010110011", -- 8882 FREE #<CONS 0 8883>
 "00000000000000000010001010110100", -- 8883 FREE #<CONS 0 8884>
 "00000000000000000010001010110101", -- 8884 FREE #<CONS 0 8885>
 "00000000000000000010001010110110", -- 8885 FREE #<CONS 0 8886>
 "00000000000000000010001010110111", -- 8886 FREE #<CONS 0 8887>
 "00000000000000000010001010111000", -- 8887 FREE #<CONS 0 8888>
 "00000000000000000010001010111001", -- 8888 FREE #<CONS 0 8889>
 "00000000000000000010001010111010", -- 8889 FREE #<CONS 0 8890>
 "00000000000000000010001010111011", -- 8890 FREE #<CONS 0 8891>
 "00000000000000000010001010111100", -- 8891 FREE #<CONS 0 8892>
 "00000000000000000010001010111101", -- 8892 FREE #<CONS 0 8893>
 "00000000000000000010001010111110", -- 8893 FREE #<CONS 0 8894>
 "00000000000000000010001010111111", -- 8894 FREE #<CONS 0 8895>
 "00000000000000000010001011000000", -- 8895 FREE #<CONS 0 8896>
 "00000000000000000010001011000001", -- 8896 FREE #<CONS 0 8897>
 "00000000000000000010001011000010", -- 8897 FREE #<CONS 0 8898>
 "00000000000000000010001011000011", -- 8898 FREE #<CONS 0 8899>
 "00000000000000000010001011000100", -- 8899 FREE #<CONS 0 8900>
 "00000000000000000010001011000101", -- 8900 FREE #<CONS 0 8901>
 "00000000000000000010001011000110", -- 8901 FREE #<CONS 0 8902>
 "00000000000000000010001011000111", -- 8902 FREE #<CONS 0 8903>
 "00000000000000000010001011001000", -- 8903 FREE #<CONS 0 8904>
 "00000000000000000010001011001001", -- 8904 FREE #<CONS 0 8905>
 "00000000000000000010001011001010", -- 8905 FREE #<CONS 0 8906>
 "00000000000000000010001011001011", -- 8906 FREE #<CONS 0 8907>
 "00000000000000000010001011001100", -- 8907 FREE #<CONS 0 8908>
 "00000000000000000010001011001101", -- 8908 FREE #<CONS 0 8909>
 "00000000000000000010001011001110", -- 8909 FREE #<CONS 0 8910>
 "00000000000000000010001011001111", -- 8910 FREE #<CONS 0 8911>
 "00000000000000000010001011010000", -- 8911 FREE #<CONS 0 8912>
 "00000000000000000010001011010001", -- 8912 FREE #<CONS 0 8913>
 "00000000000000000010001011010010", -- 8913 FREE #<CONS 0 8914>
 "00000000000000000010001011010011", -- 8914 FREE #<CONS 0 8915>
 "00000000000000000010001011010100", -- 8915 FREE #<CONS 0 8916>
 "00000000000000000010001011010101", -- 8916 FREE #<CONS 0 8917>
 "00000000000000000010001011010110", -- 8917 FREE #<CONS 0 8918>
 "00000000000000000010001011010111", -- 8918 FREE #<CONS 0 8919>
 "00000000000000000010001011011000", -- 8919 FREE #<CONS 0 8920>
 "00000000000000000010001011011001", -- 8920 FREE #<CONS 0 8921>
 "00000000000000000010001011011010", -- 8921 FREE #<CONS 0 8922>
 "00000000000000000010001011011011", -- 8922 FREE #<CONS 0 8923>
 "00000000000000000010001011011100", -- 8923 FREE #<CONS 0 8924>
 "00000000000000000010001011011101", -- 8924 FREE #<CONS 0 8925>
 "00000000000000000010001011011110", -- 8925 FREE #<CONS 0 8926>
 "00000000000000000010001011011111", -- 8926 FREE #<CONS 0 8927>
 "00000000000000000010001011100000", -- 8927 FREE #<CONS 0 8928>
 "00000000000000000010001011100001", -- 8928 FREE #<CONS 0 8929>
 "00000000000000000010001011100010", -- 8929 FREE #<CONS 0 8930>
 "00000000000000000010001011100011", -- 8930 FREE #<CONS 0 8931>
 "00000000000000000010001011100100", -- 8931 FREE #<CONS 0 8932>
 "00000000000000000010001011100101", -- 8932 FREE #<CONS 0 8933>
 "00000000000000000010001011100110", -- 8933 FREE #<CONS 0 8934>
 "00000000000000000010001011100111", -- 8934 FREE #<CONS 0 8935>
 "00000000000000000010001011101000", -- 8935 FREE #<CONS 0 8936>
 "00000000000000000010001011101001", -- 8936 FREE #<CONS 0 8937>
 "00000000000000000010001011101010", -- 8937 FREE #<CONS 0 8938>
 "00000000000000000010001011101011", -- 8938 FREE #<CONS 0 8939>
 "00000000000000000010001011101100", -- 8939 FREE #<CONS 0 8940>
 "00000000000000000010001011101101", -- 8940 FREE #<CONS 0 8941>
 "00000000000000000010001011101110", -- 8941 FREE #<CONS 0 8942>
 "00000000000000000010001011101111", -- 8942 FREE #<CONS 0 8943>
 "00000000000000000010001011110000", -- 8943 FREE #<CONS 0 8944>
 "00000000000000000010001011110001", -- 8944 FREE #<CONS 0 8945>
 "00000000000000000010001011110010", -- 8945 FREE #<CONS 0 8946>
 "00000000000000000010001011110011", -- 8946 FREE #<CONS 0 8947>
 "00000000000000000010001011110100", -- 8947 FREE #<CONS 0 8948>
 "00000000000000000010001011110101", -- 8948 FREE #<CONS 0 8949>
 "00000000000000000010001011110110", -- 8949 FREE #<CONS 0 8950>
 "00000000000000000010001011110111", -- 8950 FREE #<CONS 0 8951>
 "00000000000000000010001011111000", -- 8951 FREE #<CONS 0 8952>
 "00000000000000000010001011111001", -- 8952 FREE #<CONS 0 8953>
 "00000000000000000010001011111010", -- 8953 FREE #<CONS 0 8954>
 "00000000000000000010001011111011", -- 8954 FREE #<CONS 0 8955>
 "00000000000000000010001011111100", -- 8955 FREE #<CONS 0 8956>
 "00000000000000000010001011111101", -- 8956 FREE #<CONS 0 8957>
 "00000000000000000010001011111110", -- 8957 FREE #<CONS 0 8958>
 "00000000000000000010001011111111", -- 8958 FREE #<CONS 0 8959>
 "00000000000000000010001100000000", -- 8959 FREE #<CONS 0 8960>
 "00000000000000000010001100000001", -- 8960 FREE #<CONS 0 8961>
 "00000000000000000010001100000010", -- 8961 FREE #<CONS 0 8962>
 "00000000000000000010001100000011", -- 8962 FREE #<CONS 0 8963>
 "00000000000000000010001100000100", -- 8963 FREE #<CONS 0 8964>
 "00000000000000000010001100000101", -- 8964 FREE #<CONS 0 8965>
 "00000000000000000010001100000110", -- 8965 FREE #<CONS 0 8966>
 "00000000000000000010001100000111", -- 8966 FREE #<CONS 0 8967>
 "00000000000000000010001100001000", -- 8967 FREE #<CONS 0 8968>
 "00000000000000000010001100001001", -- 8968 FREE #<CONS 0 8969>
 "00000000000000000010001100001010", -- 8969 FREE #<CONS 0 8970>
 "00000000000000000010001100001011", -- 8970 FREE #<CONS 0 8971>
 "00000000000000000010001100001100", -- 8971 FREE #<CONS 0 8972>
 "00000000000000000010001100001101", -- 8972 FREE #<CONS 0 8973>
 "00000000000000000010001100001110", -- 8973 FREE #<CONS 0 8974>
 "00000000000000000010001100001111", -- 8974 FREE #<CONS 0 8975>
 "00000000000000000010001100010000", -- 8975 FREE #<CONS 0 8976>
 "00000000000000000010001100010001", -- 8976 FREE #<CONS 0 8977>
 "00000000000000000010001100010010", -- 8977 FREE #<CONS 0 8978>
 "00000000000000000010001100010011", -- 8978 FREE #<CONS 0 8979>
 "00000000000000000010001100010100", -- 8979 FREE #<CONS 0 8980>
 "00000000000000000010001100010101", -- 8980 FREE #<CONS 0 8981>
 "00000000000000000010001100010110", -- 8981 FREE #<CONS 0 8982>
 "00000000000000000010001100010111", -- 8982 FREE #<CONS 0 8983>
 "00000000000000000010001100011000", -- 8983 FREE #<CONS 0 8984>
 "00000000000000000010001100011001", -- 8984 FREE #<CONS 0 8985>
 "00000000000000000010001100011010", -- 8985 FREE #<CONS 0 8986>
 "00000000000000000010001100011011", -- 8986 FREE #<CONS 0 8987>
 "00000000000000000010001100011100", -- 8987 FREE #<CONS 0 8988>
 "00000000000000000010001100011101", -- 8988 FREE #<CONS 0 8989>
 "00000000000000000010001100011110", -- 8989 FREE #<CONS 0 8990>
 "00000000000000000010001100011111", -- 8990 FREE #<CONS 0 8991>
 "00000000000000000010001100100000", -- 8991 FREE #<CONS 0 8992>
 "00000000000000000010001100100001", -- 8992 FREE #<CONS 0 8993>
 "00000000000000000010001100100010", -- 8993 FREE #<CONS 0 8994>
 "00000000000000000010001100100011", -- 8994 FREE #<CONS 0 8995>
 "00000000000000000010001100100100", -- 8995 FREE #<CONS 0 8996>
 "00000000000000000010001100100101", -- 8996 FREE #<CONS 0 8997>
 "00000000000000000010001100100110", -- 8997 FREE #<CONS 0 8998>
 "00000000000000000010001100100111", -- 8998 FREE #<CONS 0 8999>
 "00000000000000000010001100101000", -- 8999 FREE #<CONS 0 9000>
 "00000000000000000010001100101001", -- 9000 FREE #<CONS 0 9001>
 "00000000000000000010001100101010", -- 9001 FREE #<CONS 0 9002>
 "00000000000000000010001100101011", -- 9002 FREE #<CONS 0 9003>
 "00000000000000000010001100101100", -- 9003 FREE #<CONS 0 9004>
 "00000000000000000010001100101101", -- 9004 FREE #<CONS 0 9005>
 "00000000000000000010001100101110", -- 9005 FREE #<CONS 0 9006>
 "00000000000000000010001100101111", -- 9006 FREE #<CONS 0 9007>
 "00000000000000000010001100110000", -- 9007 FREE #<CONS 0 9008>
 "00000000000000000010001100110001", -- 9008 FREE #<CONS 0 9009>
 "00000000000000000010001100110010", -- 9009 FREE #<CONS 0 9010>
 "00000000000000000010001100110011", -- 9010 FREE #<CONS 0 9011>
 "00000000000000000010001100110100", -- 9011 FREE #<CONS 0 9012>
 "00000000000000000010001100110101", -- 9012 FREE #<CONS 0 9013>
 "00000000000000000010001100110110", -- 9013 FREE #<CONS 0 9014>
 "00000000000000000010001100110111", -- 9014 FREE #<CONS 0 9015>
 "00000000000000000010001100111000", -- 9015 FREE #<CONS 0 9016>
 "00000000000000000010001100111001", -- 9016 FREE #<CONS 0 9017>
 "00000000000000000010001100111010", -- 9017 FREE #<CONS 0 9018>
 "00000000000000000010001100111011", -- 9018 FREE #<CONS 0 9019>
 "00000000000000000010001100111100", -- 9019 FREE #<CONS 0 9020>
 "00000000000000000010001100111101", -- 9020 FREE #<CONS 0 9021>
 "00000000000000000010001100111110", -- 9021 FREE #<CONS 0 9022>
 "00000000000000000010001100111111", -- 9022 FREE #<CONS 0 9023>
 "00000000000000000010001101000000", -- 9023 FREE #<CONS 0 9024>
 "00000000000000000010001101000001", -- 9024 FREE #<CONS 0 9025>
 "00000000000000000010001101000010", -- 9025 FREE #<CONS 0 9026>
 "00000000000000000010001101000011", -- 9026 FREE #<CONS 0 9027>
 "00000000000000000010001101000100", -- 9027 FREE #<CONS 0 9028>
 "00000000000000000010001101000101", -- 9028 FREE #<CONS 0 9029>
 "00000000000000000010001101000110", -- 9029 FREE #<CONS 0 9030>
 "00000000000000000010001101000111", -- 9030 FREE #<CONS 0 9031>
 "00000000000000000010001101001000", -- 9031 FREE #<CONS 0 9032>
 "00000000000000000010001101001001", -- 9032 FREE #<CONS 0 9033>
 "00000000000000000010001101001010", -- 9033 FREE #<CONS 0 9034>
 "00000000000000000010001101001011", -- 9034 FREE #<CONS 0 9035>
 "00000000000000000010001101001100", -- 9035 FREE #<CONS 0 9036>
 "00000000000000000010001101001101", -- 9036 FREE #<CONS 0 9037>
 "00000000000000000010001101001110", -- 9037 FREE #<CONS 0 9038>
 "00000000000000000010001101001111", -- 9038 FREE #<CONS 0 9039>
 "00000000000000000010001101010000", -- 9039 FREE #<CONS 0 9040>
 "00000000000000000010001101010001", -- 9040 FREE #<CONS 0 9041>
 "00000000000000000010001101010010", -- 9041 FREE #<CONS 0 9042>
 "00000000000000000010001101010011", -- 9042 FREE #<CONS 0 9043>
 "00000000000000000010001101010100", -- 9043 FREE #<CONS 0 9044>
 "00000000000000000010001101010101", -- 9044 FREE #<CONS 0 9045>
 "00000000000000000010001101010110", -- 9045 FREE #<CONS 0 9046>
 "00000000000000000010001101010111", -- 9046 FREE #<CONS 0 9047>
 "00000000000000000010001101011000", -- 9047 FREE #<CONS 0 9048>
 "00000000000000000010001101011001", -- 9048 FREE #<CONS 0 9049>
 "00000000000000000010001101011010", -- 9049 FREE #<CONS 0 9050>
 "00000000000000000010001101011011", -- 9050 FREE #<CONS 0 9051>
 "00000000000000000010001101011100", -- 9051 FREE #<CONS 0 9052>
 "00000000000000000010001101011101", -- 9052 FREE #<CONS 0 9053>
 "00000000000000000010001101011110", -- 9053 FREE #<CONS 0 9054>
 "00000000000000000010001101011111", -- 9054 FREE #<CONS 0 9055>
 "00000000000000000010001101100000", -- 9055 FREE #<CONS 0 9056>
 "00000000000000000010001101100001", -- 9056 FREE #<CONS 0 9057>
 "00000000000000000010001101100010", -- 9057 FREE #<CONS 0 9058>
 "00000000000000000010001101100011", -- 9058 FREE #<CONS 0 9059>
 "00000000000000000010001101100100", -- 9059 FREE #<CONS 0 9060>
 "00000000000000000010001101100101", -- 9060 FREE #<CONS 0 9061>
 "00000000000000000010001101100110", -- 9061 FREE #<CONS 0 9062>
 "00000000000000000010001101100111", -- 9062 FREE #<CONS 0 9063>
 "00000000000000000010001101101000", -- 9063 FREE #<CONS 0 9064>
 "00000000000000000010001101101001", -- 9064 FREE #<CONS 0 9065>
 "00000000000000000010001101101010", -- 9065 FREE #<CONS 0 9066>
 "00000000000000000010001101101011", -- 9066 FREE #<CONS 0 9067>
 "00000000000000000010001101101100", -- 9067 FREE #<CONS 0 9068>
 "00000000000000000010001101101101", -- 9068 FREE #<CONS 0 9069>
 "00000000000000000010001101101110", -- 9069 FREE #<CONS 0 9070>
 "00000000000000000010001101101111", -- 9070 FREE #<CONS 0 9071>
 "00000000000000000010001101110000", -- 9071 FREE #<CONS 0 9072>
 "00000000000000000010001101110001", -- 9072 FREE #<CONS 0 9073>
 "00000000000000000010001101110010", -- 9073 FREE #<CONS 0 9074>
 "00000000000000000010001101110011", -- 9074 FREE #<CONS 0 9075>
 "00000000000000000010001101110100", -- 9075 FREE #<CONS 0 9076>
 "00000000000000000010001101110101", -- 9076 FREE #<CONS 0 9077>
 "00000000000000000010001101110110", -- 9077 FREE #<CONS 0 9078>
 "00000000000000000010001101110111", -- 9078 FREE #<CONS 0 9079>
 "00000000000000000010001101111000", -- 9079 FREE #<CONS 0 9080>
 "00000000000000000010001101111001", -- 9080 FREE #<CONS 0 9081>
 "00000000000000000010001101111010", -- 9081 FREE #<CONS 0 9082>
 "00000000000000000010001101111011", -- 9082 FREE #<CONS 0 9083>
 "00000000000000000010001101111100", -- 9083 FREE #<CONS 0 9084>
 "00000000000000000010001101111101", -- 9084 FREE #<CONS 0 9085>
 "00000000000000000010001101111110", -- 9085 FREE #<CONS 0 9086>
 "00000000000000000010001101111111", -- 9086 FREE #<CONS 0 9087>
 "00000000000000000010001110000000", -- 9087 FREE #<CONS 0 9088>
 "00000000000000000010001110000001", -- 9088 FREE #<CONS 0 9089>
 "00000000000000000010001110000010", -- 9089 FREE #<CONS 0 9090>
 "00000000000000000010001110000011", -- 9090 FREE #<CONS 0 9091>
 "00000000000000000010001110000100", -- 9091 FREE #<CONS 0 9092>
 "00000000000000000010001110000101", -- 9092 FREE #<CONS 0 9093>
 "00000000000000000010001110000110", -- 9093 FREE #<CONS 0 9094>
 "00000000000000000010001110000111", -- 9094 FREE #<CONS 0 9095>
 "00000000000000000010001110001000", -- 9095 FREE #<CONS 0 9096>
 "00000000000000000010001110001001", -- 9096 FREE #<CONS 0 9097>
 "00000000000000000010001110001010", -- 9097 FREE #<CONS 0 9098>
 "00000000000000000010001110001011", -- 9098 FREE #<CONS 0 9099>
 "00000000000000000010001110001100", -- 9099 FREE #<CONS 0 9100>
 "00000000000000000010001110001101", -- 9100 FREE #<CONS 0 9101>
 "00000000000000000010001110001110", -- 9101 FREE #<CONS 0 9102>
 "00000000000000000010001110001111", -- 9102 FREE #<CONS 0 9103>
 "00000000000000000010001110010000", -- 9103 FREE #<CONS 0 9104>
 "00000000000000000010001110010001", -- 9104 FREE #<CONS 0 9105>
 "00000000000000000010001110010010", -- 9105 FREE #<CONS 0 9106>
 "00000000000000000010001110010011", -- 9106 FREE #<CONS 0 9107>
 "00000000000000000010001110010100", -- 9107 FREE #<CONS 0 9108>
 "00000000000000000010001110010101", -- 9108 FREE #<CONS 0 9109>
 "00000000000000000010001110010110", -- 9109 FREE #<CONS 0 9110>
 "00000000000000000010001110010111", -- 9110 FREE #<CONS 0 9111>
 "00000000000000000010001110011000", -- 9111 FREE #<CONS 0 9112>
 "00000000000000000010001110011001", -- 9112 FREE #<CONS 0 9113>
 "00000000000000000010001110011010", -- 9113 FREE #<CONS 0 9114>
 "00000000000000000010001110011011", -- 9114 FREE #<CONS 0 9115>
 "00000000000000000010001110011100", -- 9115 FREE #<CONS 0 9116>
 "00000000000000000010001110011101", -- 9116 FREE #<CONS 0 9117>
 "00000000000000000010001110011110", -- 9117 FREE #<CONS 0 9118>
 "00000000000000000010001110011111", -- 9118 FREE #<CONS 0 9119>
 "00000000000000000010001110100000", -- 9119 FREE #<CONS 0 9120>
 "00000000000000000010001110100001", -- 9120 FREE #<CONS 0 9121>
 "00000000000000000010001110100010", -- 9121 FREE #<CONS 0 9122>
 "00000000000000000010001110100011", -- 9122 FREE #<CONS 0 9123>
 "00000000000000000010001110100100", -- 9123 FREE #<CONS 0 9124>
 "00000000000000000010001110100101", -- 9124 FREE #<CONS 0 9125>
 "00000000000000000010001110100110", -- 9125 FREE #<CONS 0 9126>
 "00000000000000000010001110100111", -- 9126 FREE #<CONS 0 9127>
 "00000000000000000010001110101000", -- 9127 FREE #<CONS 0 9128>
 "00000000000000000010001110101001", -- 9128 FREE #<CONS 0 9129>
 "00000000000000000010001110101010", -- 9129 FREE #<CONS 0 9130>
 "00000000000000000010001110101011", -- 9130 FREE #<CONS 0 9131>
 "00000000000000000010001110101100", -- 9131 FREE #<CONS 0 9132>
 "00000000000000000010001110101101", -- 9132 FREE #<CONS 0 9133>
 "00000000000000000010001110101110", -- 9133 FREE #<CONS 0 9134>
 "00000000000000000010001110101111", -- 9134 FREE #<CONS 0 9135>
 "00000000000000000010001110110000", -- 9135 FREE #<CONS 0 9136>
 "00000000000000000010001110110001", -- 9136 FREE #<CONS 0 9137>
 "00000000000000000010001110110010", -- 9137 FREE #<CONS 0 9138>
 "00000000000000000010001110110011", -- 9138 FREE #<CONS 0 9139>
 "00000000000000000010001110110100", -- 9139 FREE #<CONS 0 9140>
 "00000000000000000010001110110101", -- 9140 FREE #<CONS 0 9141>
 "00000000000000000010001110110110", -- 9141 FREE #<CONS 0 9142>
 "00000000000000000010001110110111", -- 9142 FREE #<CONS 0 9143>
 "00000000000000000010001110111000", -- 9143 FREE #<CONS 0 9144>
 "00000000000000000010001110111001", -- 9144 FREE #<CONS 0 9145>
 "00000000000000000010001110111010", -- 9145 FREE #<CONS 0 9146>
 "00000000000000000010001110111011", -- 9146 FREE #<CONS 0 9147>
 "00000000000000000010001110111100", -- 9147 FREE #<CONS 0 9148>
 "00000000000000000010001110111101", -- 9148 FREE #<CONS 0 9149>
 "00000000000000000010001110111110", -- 9149 FREE #<CONS 0 9150>
 "00000000000000000010001110111111", -- 9150 FREE #<CONS 0 9151>
 "00000000000000000010001111000000", -- 9151 FREE #<CONS 0 9152>
 "00000000000000000010001111000001", -- 9152 FREE #<CONS 0 9153>
 "00000000000000000010001111000010", -- 9153 FREE #<CONS 0 9154>
 "00000000000000000010001111000011", -- 9154 FREE #<CONS 0 9155>
 "00000000000000000010001111000100", -- 9155 FREE #<CONS 0 9156>
 "00000000000000000010001111000101", -- 9156 FREE #<CONS 0 9157>
 "00000000000000000010001111000110", -- 9157 FREE #<CONS 0 9158>
 "00000000000000000010001111000111", -- 9158 FREE #<CONS 0 9159>
 "00000000000000000010001111001000", -- 9159 FREE #<CONS 0 9160>
 "00000000000000000010001111001001", -- 9160 FREE #<CONS 0 9161>
 "00000000000000000010001111001010", -- 9161 FREE #<CONS 0 9162>
 "00000000000000000010001111001011", -- 9162 FREE #<CONS 0 9163>
 "00000000000000000010001111001100", -- 9163 FREE #<CONS 0 9164>
 "00000000000000000010001111001101", -- 9164 FREE #<CONS 0 9165>
 "00000000000000000010001111001110", -- 9165 FREE #<CONS 0 9166>
 "00000000000000000010001111001111", -- 9166 FREE #<CONS 0 9167>
 "00000000000000000010001111010000", -- 9167 FREE #<CONS 0 9168>
 "00000000000000000010001111010001", -- 9168 FREE #<CONS 0 9169>
 "00000000000000000010001111010010", -- 9169 FREE #<CONS 0 9170>
 "00000000000000000010001111010011", -- 9170 FREE #<CONS 0 9171>
 "00000000000000000010001111010100", -- 9171 FREE #<CONS 0 9172>
 "00000000000000000010001111010101", -- 9172 FREE #<CONS 0 9173>
 "00000000000000000010001111010110", -- 9173 FREE #<CONS 0 9174>
 "00000000000000000010001111010111", -- 9174 FREE #<CONS 0 9175>
 "00000000000000000010001111011000", -- 9175 FREE #<CONS 0 9176>
 "00000000000000000010001111011001", -- 9176 FREE #<CONS 0 9177>
 "00000000000000000010001111011010", -- 9177 FREE #<CONS 0 9178>
 "00000000000000000010001111011011", -- 9178 FREE #<CONS 0 9179>
 "00000000000000000010001111011100", -- 9179 FREE #<CONS 0 9180>
 "00000000000000000010001111011101", -- 9180 FREE #<CONS 0 9181>
 "00000000000000000010001111011110", -- 9181 FREE #<CONS 0 9182>
 "00000000000000000010001111011111", -- 9182 FREE #<CONS 0 9183>
 "00000000000000000010001111100000", -- 9183 FREE #<CONS 0 9184>
 "00000000000000000010001111100001", -- 9184 FREE #<CONS 0 9185>
 "00000000000000000010001111100010", -- 9185 FREE #<CONS 0 9186>
 "00000000000000000010001111100011", -- 9186 FREE #<CONS 0 9187>
 "00000000000000000010001111100100", -- 9187 FREE #<CONS 0 9188>
 "00000000000000000010001111100101", -- 9188 FREE #<CONS 0 9189>
 "00000000000000000010001111100110", -- 9189 FREE #<CONS 0 9190>
 "00000000000000000010001111100111", -- 9190 FREE #<CONS 0 9191>
 "00000000000000000010001111101000", -- 9191 FREE #<CONS 0 9192>
 "00000000000000000010001111101001", -- 9192 FREE #<CONS 0 9193>
 "00000000000000000010001111101010", -- 9193 FREE #<CONS 0 9194>
 "00000000000000000010001111101011", -- 9194 FREE #<CONS 0 9195>
 "00000000000000000010001111101100", -- 9195 FREE #<CONS 0 9196>
 "00000000000000000010001111101101", -- 9196 FREE #<CONS 0 9197>
 "00000000000000000010001111101110", -- 9197 FREE #<CONS 0 9198>
 "00000000000000000010001111101111", -- 9198 FREE #<CONS 0 9199>
 "00000000000000000010001111110000", -- 9199 FREE #<CONS 0 9200>
 "00000000000000000010001111110001", -- 9200 FREE #<CONS 0 9201>
 "00000000000000000010001111110010", -- 9201 FREE #<CONS 0 9202>
 "00000000000000000010001111110011", -- 9202 FREE #<CONS 0 9203>
 "00000000000000000010001111110100", -- 9203 FREE #<CONS 0 9204>
 "00000000000000000010001111110101", -- 9204 FREE #<CONS 0 9205>
 "00000000000000000010001111110110", -- 9205 FREE #<CONS 0 9206>
 "00000000000000000010001111110111", -- 9206 FREE #<CONS 0 9207>
 "00000000000000000010001111111000", -- 9207 FREE #<CONS 0 9208>
 "00000000000000000010001111111001", -- 9208 FREE #<CONS 0 9209>
 "00000000000000000010001111111010", -- 9209 FREE #<CONS 0 9210>
 "00000000000000000010001111111011", -- 9210 FREE #<CONS 0 9211>
 "00000000000000000010001111111100", -- 9211 FREE #<CONS 0 9212>
 "00000000000000000010001111111101", -- 9212 FREE #<CONS 0 9213>
 "00000000000000000010001111111110", -- 9213 FREE #<CONS 0 9214>
 "00000000000000000010001111111111", -- 9214 FREE #<CONS 0 9215>
 "00000000000000000010010000000000", -- 9215 FREE #<CONS 0 9216>
 "00000000000000000010010000000001", -- 9216 FREE #<CONS 0 9217>
 "00000000000000000010010000000010", -- 9217 FREE #<CONS 0 9218>
 "00000000000000000010010000000011", -- 9218 FREE #<CONS 0 9219>
 "00000000000000000010010000000100", -- 9219 FREE #<CONS 0 9220>
 "00000000000000000010010000000101", -- 9220 FREE #<CONS 0 9221>
 "00000000000000000010010000000110", -- 9221 FREE #<CONS 0 9222>
 "00000000000000000010010000000111", -- 9222 FREE #<CONS 0 9223>
 "00000000000000000010010000001000", -- 9223 FREE #<CONS 0 9224>
 "00000000000000000010010000001001", -- 9224 FREE #<CONS 0 9225>
 "00000000000000000010010000001010", -- 9225 FREE #<CONS 0 9226>
 "00000000000000000010010000001011", -- 9226 FREE #<CONS 0 9227>
 "00000000000000000010010000001100", -- 9227 FREE #<CONS 0 9228>
 "00000000000000000010010000001101", -- 9228 FREE #<CONS 0 9229>
 "00000000000000000010010000001110", -- 9229 FREE #<CONS 0 9230>
 "00000000000000000010010000001111", -- 9230 FREE #<CONS 0 9231>
 "00000000000000000010010000010000", -- 9231 FREE #<CONS 0 9232>
 "00000000000000000010010000010001", -- 9232 FREE #<CONS 0 9233>
 "00000000000000000010010000010010", -- 9233 FREE #<CONS 0 9234>
 "00000000000000000010010000010011", -- 9234 FREE #<CONS 0 9235>
 "00000000000000000010010000010100", -- 9235 FREE #<CONS 0 9236>
 "00000000000000000010010000010101", -- 9236 FREE #<CONS 0 9237>
 "00000000000000000010010000010110", -- 9237 FREE #<CONS 0 9238>
 "00000000000000000010010000010111", -- 9238 FREE #<CONS 0 9239>
 "00000000000000000010010000011000", -- 9239 FREE #<CONS 0 9240>
 "00000000000000000010010000011001", -- 9240 FREE #<CONS 0 9241>
 "00000000000000000010010000011010", -- 9241 FREE #<CONS 0 9242>
 "00000000000000000010010000011011", -- 9242 FREE #<CONS 0 9243>
 "00000000000000000010010000011100", -- 9243 FREE #<CONS 0 9244>
 "00000000000000000010010000011101", -- 9244 FREE #<CONS 0 9245>
 "00000000000000000010010000011110", -- 9245 FREE #<CONS 0 9246>
 "00000000000000000010010000011111", -- 9246 FREE #<CONS 0 9247>
 "00000000000000000010010000100000", -- 9247 FREE #<CONS 0 9248>
 "00000000000000000010010000100001", -- 9248 FREE #<CONS 0 9249>
 "00000000000000000010010000100010", -- 9249 FREE #<CONS 0 9250>
 "00000000000000000010010000100011", -- 9250 FREE #<CONS 0 9251>
 "00000000000000000010010000100100", -- 9251 FREE #<CONS 0 9252>
 "00000000000000000010010000100101", -- 9252 FREE #<CONS 0 9253>
 "00000000000000000010010000100110", -- 9253 FREE #<CONS 0 9254>
 "00000000000000000010010000100111", -- 9254 FREE #<CONS 0 9255>
 "00000000000000000010010000101000", -- 9255 FREE #<CONS 0 9256>
 "00000000000000000010010000101001", -- 9256 FREE #<CONS 0 9257>
 "00000000000000000010010000101010", -- 9257 FREE #<CONS 0 9258>
 "00000000000000000010010000101011", -- 9258 FREE #<CONS 0 9259>
 "00000000000000000010010000101100", -- 9259 FREE #<CONS 0 9260>
 "00000000000000000010010000101101", -- 9260 FREE #<CONS 0 9261>
 "00000000000000000010010000101110", -- 9261 FREE #<CONS 0 9262>
 "00000000000000000010010000101111", -- 9262 FREE #<CONS 0 9263>
 "00000000000000000010010000110000", -- 9263 FREE #<CONS 0 9264>
 "00000000000000000010010000110001", -- 9264 FREE #<CONS 0 9265>
 "00000000000000000010010000110010", -- 9265 FREE #<CONS 0 9266>
 "00000000000000000010010000110011", -- 9266 FREE #<CONS 0 9267>
 "00000000000000000010010000110100", -- 9267 FREE #<CONS 0 9268>
 "00000000000000000010010000110101", -- 9268 FREE #<CONS 0 9269>
 "00000000000000000010010000110110", -- 9269 FREE #<CONS 0 9270>
 "00000000000000000010010000110111", -- 9270 FREE #<CONS 0 9271>
 "00000000000000000010010000111000", -- 9271 FREE #<CONS 0 9272>
 "00000000000000000010010000111001", -- 9272 FREE #<CONS 0 9273>
 "00000000000000000010010000111010", -- 9273 FREE #<CONS 0 9274>
 "00000000000000000010010000111011", -- 9274 FREE #<CONS 0 9275>
 "00000000000000000010010000111100", -- 9275 FREE #<CONS 0 9276>
 "00000000000000000010010000111101", -- 9276 FREE #<CONS 0 9277>
 "00000000000000000010010000111110", -- 9277 FREE #<CONS 0 9278>
 "00000000000000000010010000111111", -- 9278 FREE #<CONS 0 9279>
 "00000000000000000010010001000000", -- 9279 FREE #<CONS 0 9280>
 "00000000000000000010010001000001", -- 9280 FREE #<CONS 0 9281>
 "00000000000000000010010001000010", -- 9281 FREE #<CONS 0 9282>
 "00000000000000000010010001000011", -- 9282 FREE #<CONS 0 9283>
 "00000000000000000010010001000100", -- 9283 FREE #<CONS 0 9284>
 "00000000000000000010010001000101", -- 9284 FREE #<CONS 0 9285>
 "00000000000000000010010001000110", -- 9285 FREE #<CONS 0 9286>
 "00000000000000000010010001000111", -- 9286 FREE #<CONS 0 9287>
 "00000000000000000010010001001000", -- 9287 FREE #<CONS 0 9288>
 "00000000000000000010010001001001", -- 9288 FREE #<CONS 0 9289>
 "00000000000000000010010001001010", -- 9289 FREE #<CONS 0 9290>
 "00000000000000000010010001001011", -- 9290 FREE #<CONS 0 9291>
 "00000000000000000010010001001100", -- 9291 FREE #<CONS 0 9292>
 "00000000000000000010010001001101", -- 9292 FREE #<CONS 0 9293>
 "00000000000000000010010001001110", -- 9293 FREE #<CONS 0 9294>
 "00000000000000000010010001001111", -- 9294 FREE #<CONS 0 9295>
 "00000000000000000010010001010000", -- 9295 FREE #<CONS 0 9296>
 "00000000000000000010010001010001", -- 9296 FREE #<CONS 0 9297>
 "00000000000000000010010001010010", -- 9297 FREE #<CONS 0 9298>
 "00000000000000000010010001010011", -- 9298 FREE #<CONS 0 9299>
 "00000000000000000010010001010100", -- 9299 FREE #<CONS 0 9300>
 "00000000000000000010010001010101", -- 9300 FREE #<CONS 0 9301>
 "00000000000000000010010001010110", -- 9301 FREE #<CONS 0 9302>
 "00000000000000000010010001010111", -- 9302 FREE #<CONS 0 9303>
 "00000000000000000010010001011000", -- 9303 FREE #<CONS 0 9304>
 "00000000000000000010010001011001", -- 9304 FREE #<CONS 0 9305>
 "00000000000000000010010001011010", -- 9305 FREE #<CONS 0 9306>
 "00000000000000000010010001011011", -- 9306 FREE #<CONS 0 9307>
 "00000000000000000010010001011100", -- 9307 FREE #<CONS 0 9308>
 "00000000000000000010010001011101", -- 9308 FREE #<CONS 0 9309>
 "00000000000000000010010001011110", -- 9309 FREE #<CONS 0 9310>
 "00000000000000000010010001011111", -- 9310 FREE #<CONS 0 9311>
 "00000000000000000010010001100000", -- 9311 FREE #<CONS 0 9312>
 "00000000000000000010010001100001", -- 9312 FREE #<CONS 0 9313>
 "00000000000000000010010001100010", -- 9313 FREE #<CONS 0 9314>
 "00000000000000000010010001100011", -- 9314 FREE #<CONS 0 9315>
 "00000000000000000010010001100100", -- 9315 FREE #<CONS 0 9316>
 "00000000000000000010010001100101", -- 9316 FREE #<CONS 0 9317>
 "00000000000000000010010001100110", -- 9317 FREE #<CONS 0 9318>
 "00000000000000000010010001100111", -- 9318 FREE #<CONS 0 9319>
 "00000000000000000010010001101000", -- 9319 FREE #<CONS 0 9320>
 "00000000000000000010010001101001", -- 9320 FREE #<CONS 0 9321>
 "00000000000000000010010001101010", -- 9321 FREE #<CONS 0 9322>
 "00000000000000000010010001101011", -- 9322 FREE #<CONS 0 9323>
 "00000000000000000010010001101100", -- 9323 FREE #<CONS 0 9324>
 "00000000000000000010010001101101", -- 9324 FREE #<CONS 0 9325>
 "00000000000000000010010001101110", -- 9325 FREE #<CONS 0 9326>
 "00000000000000000010010001101111", -- 9326 FREE #<CONS 0 9327>
 "00000000000000000010010001110000", -- 9327 FREE #<CONS 0 9328>
 "00000000000000000010010001110001", -- 9328 FREE #<CONS 0 9329>
 "00000000000000000010010001110010", -- 9329 FREE #<CONS 0 9330>
 "00000000000000000010010001110011", -- 9330 FREE #<CONS 0 9331>
 "00000000000000000010010001110100", -- 9331 FREE #<CONS 0 9332>
 "00000000000000000010010001110101", -- 9332 FREE #<CONS 0 9333>
 "00000000000000000010010001110110", -- 9333 FREE #<CONS 0 9334>
 "00000000000000000010010001110111", -- 9334 FREE #<CONS 0 9335>
 "00000000000000000010010001111000", -- 9335 FREE #<CONS 0 9336>
 "00000000000000000010010001111001", -- 9336 FREE #<CONS 0 9337>
 "00000000000000000010010001111010", -- 9337 FREE #<CONS 0 9338>
 "00000000000000000010010001111011", -- 9338 FREE #<CONS 0 9339>
 "00000000000000000010010001111100", -- 9339 FREE #<CONS 0 9340>
 "00000000000000000010010001111101", -- 9340 FREE #<CONS 0 9341>
 "00000000000000000010010001111110", -- 9341 FREE #<CONS 0 9342>
 "00000000000000000010010001111111", -- 9342 FREE #<CONS 0 9343>
 "00000000000000000010010010000000", -- 9343 FREE #<CONS 0 9344>
 "00000000000000000010010010000001", -- 9344 FREE #<CONS 0 9345>
 "00000000000000000010010010000010", -- 9345 FREE #<CONS 0 9346>
 "00000000000000000010010010000011", -- 9346 FREE #<CONS 0 9347>
 "00000000000000000010010010000100", -- 9347 FREE #<CONS 0 9348>
 "00000000000000000010010010000101", -- 9348 FREE #<CONS 0 9349>
 "00000000000000000010010010000110", -- 9349 FREE #<CONS 0 9350>
 "00000000000000000010010010000111", -- 9350 FREE #<CONS 0 9351>
 "00000000000000000010010010001000", -- 9351 FREE #<CONS 0 9352>
 "00000000000000000010010010001001", -- 9352 FREE #<CONS 0 9353>
 "00000000000000000010010010001010", -- 9353 FREE #<CONS 0 9354>
 "00000000000000000010010010001011", -- 9354 FREE #<CONS 0 9355>
 "00000000000000000010010010001100", -- 9355 FREE #<CONS 0 9356>
 "00000000000000000010010010001101", -- 9356 FREE #<CONS 0 9357>
 "00000000000000000010010010001110", -- 9357 FREE #<CONS 0 9358>
 "00000000000000000010010010001111", -- 9358 FREE #<CONS 0 9359>
 "00000000000000000010010010010000", -- 9359 FREE #<CONS 0 9360>
 "00000000000000000010010010010001", -- 9360 FREE #<CONS 0 9361>
 "00000000000000000010010010010010", -- 9361 FREE #<CONS 0 9362>
 "00000000000000000010010010010011", -- 9362 FREE #<CONS 0 9363>
 "00000000000000000010010010010100", -- 9363 FREE #<CONS 0 9364>
 "00000000000000000010010010010101", -- 9364 FREE #<CONS 0 9365>
 "00000000000000000010010010010110", -- 9365 FREE #<CONS 0 9366>
 "00000000000000000010010010010111", -- 9366 FREE #<CONS 0 9367>
 "00000000000000000010010010011000", -- 9367 FREE #<CONS 0 9368>
 "00000000000000000010010010011001", -- 9368 FREE #<CONS 0 9369>
 "00000000000000000010010010011010", -- 9369 FREE #<CONS 0 9370>
 "00000000000000000010010010011011", -- 9370 FREE #<CONS 0 9371>
 "00000000000000000010010010011100", -- 9371 FREE #<CONS 0 9372>
 "00000000000000000010010010011101", -- 9372 FREE #<CONS 0 9373>
 "00000000000000000010010010011110", -- 9373 FREE #<CONS 0 9374>
 "00000000000000000010010010011111", -- 9374 FREE #<CONS 0 9375>
 "00000000000000000010010010100000", -- 9375 FREE #<CONS 0 9376>
 "00000000000000000010010010100001", -- 9376 FREE #<CONS 0 9377>
 "00000000000000000010010010100010", -- 9377 FREE #<CONS 0 9378>
 "00000000000000000010010010100011", -- 9378 FREE #<CONS 0 9379>
 "00000000000000000010010010100100", -- 9379 FREE #<CONS 0 9380>
 "00000000000000000010010010100101", -- 9380 FREE #<CONS 0 9381>
 "00000000000000000010010010100110", -- 9381 FREE #<CONS 0 9382>
 "00000000000000000010010010100111", -- 9382 FREE #<CONS 0 9383>
 "00000000000000000010010010101000", -- 9383 FREE #<CONS 0 9384>
 "00000000000000000010010010101001", -- 9384 FREE #<CONS 0 9385>
 "00000000000000000010010010101010", -- 9385 FREE #<CONS 0 9386>
 "00000000000000000010010010101011", -- 9386 FREE #<CONS 0 9387>
 "00000000000000000010010010101100", -- 9387 FREE #<CONS 0 9388>
 "00000000000000000010010010101101", -- 9388 FREE #<CONS 0 9389>
 "00000000000000000010010010101110", -- 9389 FREE #<CONS 0 9390>
 "00000000000000000010010010101111", -- 9390 FREE #<CONS 0 9391>
 "00000000000000000010010010110000", -- 9391 FREE #<CONS 0 9392>
 "00000000000000000010010010110001", -- 9392 FREE #<CONS 0 9393>
 "00000000000000000010010010110010", -- 9393 FREE #<CONS 0 9394>
 "00000000000000000010010010110011", -- 9394 FREE #<CONS 0 9395>
 "00000000000000000010010010110100", -- 9395 FREE #<CONS 0 9396>
 "00000000000000000010010010110101", -- 9396 FREE #<CONS 0 9397>
 "00000000000000000010010010110110", -- 9397 FREE #<CONS 0 9398>
 "00000000000000000010010010110111", -- 9398 FREE #<CONS 0 9399>
 "00000000000000000010010010111000", -- 9399 FREE #<CONS 0 9400>
 "00000000000000000010010010111001", -- 9400 FREE #<CONS 0 9401>
 "00000000000000000010010010111010", -- 9401 FREE #<CONS 0 9402>
 "00000000000000000010010010111011", -- 9402 FREE #<CONS 0 9403>
 "00000000000000000010010010111100", -- 9403 FREE #<CONS 0 9404>
 "00000000000000000010010010111101", -- 9404 FREE #<CONS 0 9405>
 "00000000000000000010010010111110", -- 9405 FREE #<CONS 0 9406>
 "00000000000000000010010010111111", -- 9406 FREE #<CONS 0 9407>
 "00000000000000000010010011000000", -- 9407 FREE #<CONS 0 9408>
 "00000000000000000010010011000001", -- 9408 FREE #<CONS 0 9409>
 "00000000000000000010010011000010", -- 9409 FREE #<CONS 0 9410>
 "00000000000000000010010011000011", -- 9410 FREE #<CONS 0 9411>
 "00000000000000000010010011000100", -- 9411 FREE #<CONS 0 9412>
 "00000000000000000010010011000101", -- 9412 FREE #<CONS 0 9413>
 "00000000000000000010010011000110", -- 9413 FREE #<CONS 0 9414>
 "00000000000000000010010011000111", -- 9414 FREE #<CONS 0 9415>
 "00000000000000000010010011001000", -- 9415 FREE #<CONS 0 9416>
 "00000000000000000010010011001001", -- 9416 FREE #<CONS 0 9417>
 "00000000000000000010010011001010", -- 9417 FREE #<CONS 0 9418>
 "00000000000000000010010011001011", -- 9418 FREE #<CONS 0 9419>
 "00000000000000000010010011001100", -- 9419 FREE #<CONS 0 9420>
 "00000000000000000010010011001101", -- 9420 FREE #<CONS 0 9421>
 "00000000000000000010010011001110", -- 9421 FREE #<CONS 0 9422>
 "00000000000000000010010011001111", -- 9422 FREE #<CONS 0 9423>
 "00000000000000000010010011010000", -- 9423 FREE #<CONS 0 9424>
 "00000000000000000010010011010001", -- 9424 FREE #<CONS 0 9425>
 "00000000000000000010010011010010", -- 9425 FREE #<CONS 0 9426>
 "00000000000000000010010011010011", -- 9426 FREE #<CONS 0 9427>
 "00000000000000000010010011010100", -- 9427 FREE #<CONS 0 9428>
 "00000000000000000010010011010101", -- 9428 FREE #<CONS 0 9429>
 "00000000000000000010010011010110", -- 9429 FREE #<CONS 0 9430>
 "00000000000000000010010011010111", -- 9430 FREE #<CONS 0 9431>
 "00000000000000000010010011011000", -- 9431 FREE #<CONS 0 9432>
 "00000000000000000010010011011001", -- 9432 FREE #<CONS 0 9433>
 "00000000000000000010010011011010", -- 9433 FREE #<CONS 0 9434>
 "00000000000000000010010011011011", -- 9434 FREE #<CONS 0 9435>
 "00000000000000000010010011011100", -- 9435 FREE #<CONS 0 9436>
 "00000000000000000010010011011101", -- 9436 FREE #<CONS 0 9437>
 "00000000000000000010010011011110", -- 9437 FREE #<CONS 0 9438>
 "00000000000000000010010011011111", -- 9438 FREE #<CONS 0 9439>
 "00000000000000000010010011100000", -- 9439 FREE #<CONS 0 9440>
 "00000000000000000010010011100001", -- 9440 FREE #<CONS 0 9441>
 "00000000000000000010010011100010", -- 9441 FREE #<CONS 0 9442>
 "00000000000000000010010011100011", -- 9442 FREE #<CONS 0 9443>
 "00000000000000000010010011100100", -- 9443 FREE #<CONS 0 9444>
 "00000000000000000010010011100101", -- 9444 FREE #<CONS 0 9445>
 "00000000000000000010010011100110", -- 9445 FREE #<CONS 0 9446>
 "00000000000000000010010011100111", -- 9446 FREE #<CONS 0 9447>
 "00000000000000000010010011101000", -- 9447 FREE #<CONS 0 9448>
 "00000000000000000010010011101001", -- 9448 FREE #<CONS 0 9449>
 "00000000000000000010010011101010", -- 9449 FREE #<CONS 0 9450>
 "00000000000000000010010011101011", -- 9450 FREE #<CONS 0 9451>
 "00000000000000000010010011101100", -- 9451 FREE #<CONS 0 9452>
 "00000000000000000010010011101101", -- 9452 FREE #<CONS 0 9453>
 "00000000000000000010010011101110", -- 9453 FREE #<CONS 0 9454>
 "00000000000000000010010011101111", -- 9454 FREE #<CONS 0 9455>
 "00000000000000000010010011110000", -- 9455 FREE #<CONS 0 9456>
 "00000000000000000010010011110001", -- 9456 FREE #<CONS 0 9457>
 "00000000000000000010010011110010", -- 9457 FREE #<CONS 0 9458>
 "00000000000000000010010011110011", -- 9458 FREE #<CONS 0 9459>
 "00000000000000000010010011110100", -- 9459 FREE #<CONS 0 9460>
 "00000000000000000010010011110101", -- 9460 FREE #<CONS 0 9461>
 "00000000000000000010010011110110", -- 9461 FREE #<CONS 0 9462>
 "00000000000000000010010011110111", -- 9462 FREE #<CONS 0 9463>
 "00000000000000000010010011111000", -- 9463 FREE #<CONS 0 9464>
 "00000000000000000010010011111001", -- 9464 FREE #<CONS 0 9465>
 "00000000000000000010010011111010", -- 9465 FREE #<CONS 0 9466>
 "00000000000000000010010011111011", -- 9466 FREE #<CONS 0 9467>
 "00000000000000000010010011111100", -- 9467 FREE #<CONS 0 9468>
 "00000000000000000010010011111101", -- 9468 FREE #<CONS 0 9469>
 "00000000000000000010010011111110", -- 9469 FREE #<CONS 0 9470>
 "00000000000000000010010011111111", -- 9470 FREE #<CONS 0 9471>
 "00000000000000000010010100000000", -- 9471 FREE #<CONS 0 9472>
 "00000000000000000010010100000001", -- 9472 FREE #<CONS 0 9473>
 "00000000000000000010010100000010", -- 9473 FREE #<CONS 0 9474>
 "00000000000000000010010100000011", -- 9474 FREE #<CONS 0 9475>
 "00000000000000000010010100000100", -- 9475 FREE #<CONS 0 9476>
 "00000000000000000010010100000101", -- 9476 FREE #<CONS 0 9477>
 "00000000000000000010010100000110", -- 9477 FREE #<CONS 0 9478>
 "00000000000000000010010100000111", -- 9478 FREE #<CONS 0 9479>
 "00000000000000000010010100001000", -- 9479 FREE #<CONS 0 9480>
 "00000000000000000010010100001001", -- 9480 FREE #<CONS 0 9481>
 "00000000000000000010010100001010", -- 9481 FREE #<CONS 0 9482>
 "00000000000000000010010100001011", -- 9482 FREE #<CONS 0 9483>
 "00000000000000000010010100001100", -- 9483 FREE #<CONS 0 9484>
 "00000000000000000010010100001101", -- 9484 FREE #<CONS 0 9485>
 "00000000000000000010010100001110", -- 9485 FREE #<CONS 0 9486>
 "00000000000000000010010100001111", -- 9486 FREE #<CONS 0 9487>
 "00000000000000000010010100010000", -- 9487 FREE #<CONS 0 9488>
 "00000000000000000010010100010001", -- 9488 FREE #<CONS 0 9489>
 "00000000000000000010010100010010", -- 9489 FREE #<CONS 0 9490>
 "00000000000000000010010100010011", -- 9490 FREE #<CONS 0 9491>
 "00000000000000000010010100010100", -- 9491 FREE #<CONS 0 9492>
 "00000000000000000010010100010101", -- 9492 FREE #<CONS 0 9493>
 "00000000000000000010010100010110", -- 9493 FREE #<CONS 0 9494>
 "00000000000000000010010100010111", -- 9494 FREE #<CONS 0 9495>
 "00000000000000000010010100011000", -- 9495 FREE #<CONS 0 9496>
 "00000000000000000010010100011001", -- 9496 FREE #<CONS 0 9497>
 "00000000000000000010010100011010", -- 9497 FREE #<CONS 0 9498>
 "00000000000000000010010100011011", -- 9498 FREE #<CONS 0 9499>
 "00000000000000000010010100011100", -- 9499 FREE #<CONS 0 9500>
 "00000000000000000010010100011101", -- 9500 FREE #<CONS 0 9501>
 "00000000000000000010010100011110", -- 9501 FREE #<CONS 0 9502>
 "00000000000000000010010100011111", -- 9502 FREE #<CONS 0 9503>
 "00000000000000000010010100100000", -- 9503 FREE #<CONS 0 9504>
 "00000000000000000010010100100001", -- 9504 FREE #<CONS 0 9505>
 "00000000000000000010010100100010", -- 9505 FREE #<CONS 0 9506>
 "00000000000000000010010100100011", -- 9506 FREE #<CONS 0 9507>
 "00000000000000000010010100100100", -- 9507 FREE #<CONS 0 9508>
 "00000000000000000010010100100101", -- 9508 FREE #<CONS 0 9509>
 "00000000000000000010010100100110", -- 9509 FREE #<CONS 0 9510>
 "00000000000000000010010100100111", -- 9510 FREE #<CONS 0 9511>
 "00000000000000000010010100101000", -- 9511 FREE #<CONS 0 9512>
 "00000000000000000010010100101001", -- 9512 FREE #<CONS 0 9513>
 "00000000000000000010010100101010", -- 9513 FREE #<CONS 0 9514>
 "00000000000000000010010100101011", -- 9514 FREE #<CONS 0 9515>
 "00000000000000000010010100101100", -- 9515 FREE #<CONS 0 9516>
 "00000000000000000010010100101101", -- 9516 FREE #<CONS 0 9517>
 "00000000000000000010010100101110", -- 9517 FREE #<CONS 0 9518>
 "00000000000000000010010100101111", -- 9518 FREE #<CONS 0 9519>
 "00000000000000000010010100110000", -- 9519 FREE #<CONS 0 9520>
 "00000000000000000010010100110001", -- 9520 FREE #<CONS 0 9521>
 "00000000000000000010010100110010", -- 9521 FREE #<CONS 0 9522>
 "00000000000000000010010100110011", -- 9522 FREE #<CONS 0 9523>
 "00000000000000000010010100110100", -- 9523 FREE #<CONS 0 9524>
 "00000000000000000010010100110101", -- 9524 FREE #<CONS 0 9525>
 "00000000000000000010010100110110", -- 9525 FREE #<CONS 0 9526>
 "00000000000000000010010100110111", -- 9526 FREE #<CONS 0 9527>
 "00000000000000000010010100111000", -- 9527 FREE #<CONS 0 9528>
 "00000000000000000010010100111001", -- 9528 FREE #<CONS 0 9529>
 "00000000000000000010010100111010", -- 9529 FREE #<CONS 0 9530>
 "00000000000000000010010100111011", -- 9530 FREE #<CONS 0 9531>
 "00000000000000000010010100111100", -- 9531 FREE #<CONS 0 9532>
 "00000000000000000010010100111101", -- 9532 FREE #<CONS 0 9533>
 "00000000000000000010010100111110", -- 9533 FREE #<CONS 0 9534>
 "00000000000000000010010100111111", -- 9534 FREE #<CONS 0 9535>
 "00000000000000000010010101000000", -- 9535 FREE #<CONS 0 9536>
 "00000000000000000010010101000001", -- 9536 FREE #<CONS 0 9537>
 "00000000000000000010010101000010", -- 9537 FREE #<CONS 0 9538>
 "00000000000000000010010101000011", -- 9538 FREE #<CONS 0 9539>
 "00000000000000000010010101000100", -- 9539 FREE #<CONS 0 9540>
 "00000000000000000010010101000101", -- 9540 FREE #<CONS 0 9541>
 "00000000000000000010010101000110", -- 9541 FREE #<CONS 0 9542>
 "00000000000000000010010101000111", -- 9542 FREE #<CONS 0 9543>
 "00000000000000000010010101001000", -- 9543 FREE #<CONS 0 9544>
 "00000000000000000010010101001001", -- 9544 FREE #<CONS 0 9545>
 "00000000000000000010010101001010", -- 9545 FREE #<CONS 0 9546>
 "00000000000000000010010101001011", -- 9546 FREE #<CONS 0 9547>
 "00000000000000000010010101001100", -- 9547 FREE #<CONS 0 9548>
 "00000000000000000010010101001101", -- 9548 FREE #<CONS 0 9549>
 "00000000000000000010010101001110", -- 9549 FREE #<CONS 0 9550>
 "00000000000000000010010101001111", -- 9550 FREE #<CONS 0 9551>
 "00000000000000000010010101010000", -- 9551 FREE #<CONS 0 9552>
 "00000000000000000010010101010001", -- 9552 FREE #<CONS 0 9553>
 "00000000000000000010010101010010", -- 9553 FREE #<CONS 0 9554>
 "00000000000000000010010101010011", -- 9554 FREE #<CONS 0 9555>
 "00000000000000000010010101010100", -- 9555 FREE #<CONS 0 9556>
 "00000000000000000010010101010101", -- 9556 FREE #<CONS 0 9557>
 "00000000000000000010010101010110", -- 9557 FREE #<CONS 0 9558>
 "00000000000000000010010101010111", -- 9558 FREE #<CONS 0 9559>
 "00000000000000000010010101011000", -- 9559 FREE #<CONS 0 9560>
 "00000000000000000010010101011001", -- 9560 FREE #<CONS 0 9561>
 "00000000000000000010010101011010", -- 9561 FREE #<CONS 0 9562>
 "00000000000000000010010101011011", -- 9562 FREE #<CONS 0 9563>
 "00000000000000000010010101011100", -- 9563 FREE #<CONS 0 9564>
 "00000000000000000010010101011101", -- 9564 FREE #<CONS 0 9565>
 "00000000000000000010010101011110", -- 9565 FREE #<CONS 0 9566>
 "00000000000000000010010101011111", -- 9566 FREE #<CONS 0 9567>
 "00000000000000000010010101100000", -- 9567 FREE #<CONS 0 9568>
 "00000000000000000010010101100001", -- 9568 FREE #<CONS 0 9569>
 "00000000000000000010010101100010", -- 9569 FREE #<CONS 0 9570>
 "00000000000000000010010101100011", -- 9570 FREE #<CONS 0 9571>
 "00000000000000000010010101100100", -- 9571 FREE #<CONS 0 9572>
 "00000000000000000010010101100101", -- 9572 FREE #<CONS 0 9573>
 "00000000000000000010010101100110", -- 9573 FREE #<CONS 0 9574>
 "00000000000000000010010101100111", -- 9574 FREE #<CONS 0 9575>
 "00000000000000000010010101101000", -- 9575 FREE #<CONS 0 9576>
 "00000000000000000010010101101001", -- 9576 FREE #<CONS 0 9577>
 "00000000000000000010010101101010", -- 9577 FREE #<CONS 0 9578>
 "00000000000000000010010101101011", -- 9578 FREE #<CONS 0 9579>
 "00000000000000000010010101101100", -- 9579 FREE #<CONS 0 9580>
 "00000000000000000010010101101101", -- 9580 FREE #<CONS 0 9581>
 "00000000000000000010010101101110", -- 9581 FREE #<CONS 0 9582>
 "00000000000000000010010101101111", -- 9582 FREE #<CONS 0 9583>
 "00000000000000000010010101110000", -- 9583 FREE #<CONS 0 9584>
 "00000000000000000010010101110001", -- 9584 FREE #<CONS 0 9585>
 "00000000000000000010010101110010", -- 9585 FREE #<CONS 0 9586>
 "00000000000000000010010101110011", -- 9586 FREE #<CONS 0 9587>
 "00000000000000000010010101110100", -- 9587 FREE #<CONS 0 9588>
 "00000000000000000010010101110101", -- 9588 FREE #<CONS 0 9589>
 "00000000000000000010010101110110", -- 9589 FREE #<CONS 0 9590>
 "00000000000000000010010101110111", -- 9590 FREE #<CONS 0 9591>
 "00000000000000000010010101111000", -- 9591 FREE #<CONS 0 9592>
 "00000000000000000010010101111001", -- 9592 FREE #<CONS 0 9593>
 "00000000000000000010010101111010", -- 9593 FREE #<CONS 0 9594>
 "00000000000000000010010101111011", -- 9594 FREE #<CONS 0 9595>
 "00000000000000000010010101111100", -- 9595 FREE #<CONS 0 9596>
 "00000000000000000010010101111101", -- 9596 FREE #<CONS 0 9597>
 "00000000000000000010010101111110", -- 9597 FREE #<CONS 0 9598>
 "00000000000000000010010101111111", -- 9598 FREE #<CONS 0 9599>
 "00000000000000000010010110000000", -- 9599 FREE #<CONS 0 9600>
 "00000000000000000010010110000001", -- 9600 FREE #<CONS 0 9601>
 "00000000000000000010010110000010", -- 9601 FREE #<CONS 0 9602>
 "00000000000000000010010110000011", -- 9602 FREE #<CONS 0 9603>
 "00000000000000000010010110000100", -- 9603 FREE #<CONS 0 9604>
 "00000000000000000010010110000101", -- 9604 FREE #<CONS 0 9605>
 "00000000000000000010010110000110", -- 9605 FREE #<CONS 0 9606>
 "00000000000000000010010110000111", -- 9606 FREE #<CONS 0 9607>
 "00000000000000000010010110001000", -- 9607 FREE #<CONS 0 9608>
 "00000000000000000010010110001001", -- 9608 FREE #<CONS 0 9609>
 "00000000000000000010010110001010", -- 9609 FREE #<CONS 0 9610>
 "00000000000000000010010110001011", -- 9610 FREE #<CONS 0 9611>
 "00000000000000000010010110001100", -- 9611 FREE #<CONS 0 9612>
 "00000000000000000010010110001101", -- 9612 FREE #<CONS 0 9613>
 "00000000000000000010010110001110", -- 9613 FREE #<CONS 0 9614>
 "00000000000000000010010110001111", -- 9614 FREE #<CONS 0 9615>
 "00000000000000000010010110010000", -- 9615 FREE #<CONS 0 9616>
 "00000000000000000010010110010001", -- 9616 FREE #<CONS 0 9617>
 "00000000000000000010010110010010", -- 9617 FREE #<CONS 0 9618>
 "00000000000000000010010110010011", -- 9618 FREE #<CONS 0 9619>
 "00000000000000000010010110010100", -- 9619 FREE #<CONS 0 9620>
 "00000000000000000010010110010101", -- 9620 FREE #<CONS 0 9621>
 "00000000000000000010010110010110", -- 9621 FREE #<CONS 0 9622>
 "00000000000000000010010110010111", -- 9622 FREE #<CONS 0 9623>
 "00000000000000000010010110011000", -- 9623 FREE #<CONS 0 9624>
 "00000000000000000010010110011001", -- 9624 FREE #<CONS 0 9625>
 "00000000000000000010010110011010", -- 9625 FREE #<CONS 0 9626>
 "00000000000000000010010110011011", -- 9626 FREE #<CONS 0 9627>
 "00000000000000000010010110011100", -- 9627 FREE #<CONS 0 9628>
 "00000000000000000010010110011101", -- 9628 FREE #<CONS 0 9629>
 "00000000000000000010010110011110", -- 9629 FREE #<CONS 0 9630>
 "00000000000000000010010110011111", -- 9630 FREE #<CONS 0 9631>
 "00000000000000000010010110100000", -- 9631 FREE #<CONS 0 9632>
 "00000000000000000010010110100001", -- 9632 FREE #<CONS 0 9633>
 "00000000000000000010010110100010", -- 9633 FREE #<CONS 0 9634>
 "00000000000000000010010110100011", -- 9634 FREE #<CONS 0 9635>
 "00000000000000000010010110100100", -- 9635 FREE #<CONS 0 9636>
 "00000000000000000010010110100101", -- 9636 FREE #<CONS 0 9637>
 "00000000000000000010010110100110", -- 9637 FREE #<CONS 0 9638>
 "00000000000000000010010110100111", -- 9638 FREE #<CONS 0 9639>
 "00000000000000000010010110101000", -- 9639 FREE #<CONS 0 9640>
 "00000000000000000010010110101001", -- 9640 FREE #<CONS 0 9641>
 "00000000000000000010010110101010", -- 9641 FREE #<CONS 0 9642>
 "00000000000000000010010110101011", -- 9642 FREE #<CONS 0 9643>
 "00000000000000000010010110101100", -- 9643 FREE #<CONS 0 9644>
 "00000000000000000010010110101101", -- 9644 FREE #<CONS 0 9645>
 "00000000000000000010010110101110", -- 9645 FREE #<CONS 0 9646>
 "00000000000000000010010110101111", -- 9646 FREE #<CONS 0 9647>
 "00000000000000000010010110110000", -- 9647 FREE #<CONS 0 9648>
 "00000000000000000010010110110001", -- 9648 FREE #<CONS 0 9649>
 "00000000000000000010010110110010", -- 9649 FREE #<CONS 0 9650>
 "00000000000000000010010110110011", -- 9650 FREE #<CONS 0 9651>
 "00000000000000000010010110110100", -- 9651 FREE #<CONS 0 9652>
 "00000000000000000010010110110101", -- 9652 FREE #<CONS 0 9653>
 "00000000000000000010010110110110", -- 9653 FREE #<CONS 0 9654>
 "00000000000000000010010110110111", -- 9654 FREE #<CONS 0 9655>
 "00000000000000000010010110111000", -- 9655 FREE #<CONS 0 9656>
 "00000000000000000010010110111001", -- 9656 FREE #<CONS 0 9657>
 "00000000000000000010010110111010", -- 9657 FREE #<CONS 0 9658>
 "00000000000000000010010110111011", -- 9658 FREE #<CONS 0 9659>
 "00000000000000000010010110111100", -- 9659 FREE #<CONS 0 9660>
 "00000000000000000010010110111101", -- 9660 FREE #<CONS 0 9661>
 "00000000000000000010010110111110", -- 9661 FREE #<CONS 0 9662>
 "00000000000000000010010110111111", -- 9662 FREE #<CONS 0 9663>
 "00000000000000000010010111000000", -- 9663 FREE #<CONS 0 9664>
 "00000000000000000010010111000001", -- 9664 FREE #<CONS 0 9665>
 "00000000000000000010010111000010", -- 9665 FREE #<CONS 0 9666>
 "00000000000000000010010111000011", -- 9666 FREE #<CONS 0 9667>
 "00000000000000000010010111000100", -- 9667 FREE #<CONS 0 9668>
 "00000000000000000010010111000101", -- 9668 FREE #<CONS 0 9669>
 "00000000000000000010010111000110", -- 9669 FREE #<CONS 0 9670>
 "00000000000000000010010111000111", -- 9670 FREE #<CONS 0 9671>
 "00000000000000000010010111001000", -- 9671 FREE #<CONS 0 9672>
 "00000000000000000010010111001001", -- 9672 FREE #<CONS 0 9673>
 "00000000000000000010010111001010", -- 9673 FREE #<CONS 0 9674>
 "00000000000000000010010111001011", -- 9674 FREE #<CONS 0 9675>
 "00000000000000000010010111001100", -- 9675 FREE #<CONS 0 9676>
 "00000000000000000010010111001101", -- 9676 FREE #<CONS 0 9677>
 "00000000000000000010010111001110", -- 9677 FREE #<CONS 0 9678>
 "00000000000000000010010111001111", -- 9678 FREE #<CONS 0 9679>
 "00000000000000000010010111010000", -- 9679 FREE #<CONS 0 9680>
 "00000000000000000010010111010001", -- 9680 FREE #<CONS 0 9681>
 "00000000000000000010010111010010", -- 9681 FREE #<CONS 0 9682>
 "00000000000000000010010111010011", -- 9682 FREE #<CONS 0 9683>
 "00000000000000000010010111010100", -- 9683 FREE #<CONS 0 9684>
 "00000000000000000010010111010101", -- 9684 FREE #<CONS 0 9685>
 "00000000000000000010010111010110", -- 9685 FREE #<CONS 0 9686>
 "00000000000000000010010111010111", -- 9686 FREE #<CONS 0 9687>
 "00000000000000000010010111011000", -- 9687 FREE #<CONS 0 9688>
 "00000000000000000010010111011001", -- 9688 FREE #<CONS 0 9689>
 "00000000000000000010010111011010", -- 9689 FREE #<CONS 0 9690>
 "00000000000000000010010111011011", -- 9690 FREE #<CONS 0 9691>
 "00000000000000000010010111011100", -- 9691 FREE #<CONS 0 9692>
 "00000000000000000010010111011101", -- 9692 FREE #<CONS 0 9693>
 "00000000000000000010010111011110", -- 9693 FREE #<CONS 0 9694>
 "00000000000000000010010111011111", -- 9694 FREE #<CONS 0 9695>
 "00000000000000000010010111100000", -- 9695 FREE #<CONS 0 9696>
 "00000000000000000010010111100001", -- 9696 FREE #<CONS 0 9697>
 "00000000000000000010010111100010", -- 9697 FREE #<CONS 0 9698>
 "00000000000000000010010111100011", -- 9698 FREE #<CONS 0 9699>
 "00000000000000000010010111100100", -- 9699 FREE #<CONS 0 9700>
 "00000000000000000010010111100101", -- 9700 FREE #<CONS 0 9701>
 "00000000000000000010010111100110", -- 9701 FREE #<CONS 0 9702>
 "00000000000000000010010111100111", -- 9702 FREE #<CONS 0 9703>
 "00000000000000000010010111101000", -- 9703 FREE #<CONS 0 9704>
 "00000000000000000010010111101001", -- 9704 FREE #<CONS 0 9705>
 "00000000000000000010010111101010", -- 9705 FREE #<CONS 0 9706>
 "00000000000000000010010111101011", -- 9706 FREE #<CONS 0 9707>
 "00000000000000000010010111101100", -- 9707 FREE #<CONS 0 9708>
 "00000000000000000010010111101101", -- 9708 FREE #<CONS 0 9709>
 "00000000000000000010010111101110", -- 9709 FREE #<CONS 0 9710>
 "00000000000000000010010111101111", -- 9710 FREE #<CONS 0 9711>
 "00000000000000000010010111110000", -- 9711 FREE #<CONS 0 9712>
 "00000000000000000010010111110001", -- 9712 FREE #<CONS 0 9713>
 "00000000000000000010010111110010", -- 9713 FREE #<CONS 0 9714>
 "00000000000000000010010111110011", -- 9714 FREE #<CONS 0 9715>
 "00000000000000000010010111110100", -- 9715 FREE #<CONS 0 9716>
 "00000000000000000010010111110101", -- 9716 FREE #<CONS 0 9717>
 "00000000000000000010010111110110", -- 9717 FREE #<CONS 0 9718>
 "00000000000000000010010111110111", -- 9718 FREE #<CONS 0 9719>
 "00000000000000000010010111111000", -- 9719 FREE #<CONS 0 9720>
 "00000000000000000010010111111001", -- 9720 FREE #<CONS 0 9721>
 "00000000000000000010010111111010", -- 9721 FREE #<CONS 0 9722>
 "00000000000000000010010111111011", -- 9722 FREE #<CONS 0 9723>
 "00000000000000000010010111111100", -- 9723 FREE #<CONS 0 9724>
 "00000000000000000010010111111101", -- 9724 FREE #<CONS 0 9725>
 "00000000000000000010010111111110", -- 9725 FREE #<CONS 0 9726>
 "00000000000000000010010111111111", -- 9726 FREE #<CONS 0 9727>
 "00000000000000000010011000000000", -- 9727 FREE #<CONS 0 9728>
 "00000000000000000010011000000001", -- 9728 FREE #<CONS 0 9729>
 "00000000000000000010011000000010", -- 9729 FREE #<CONS 0 9730>
 "00000000000000000010011000000011", -- 9730 FREE #<CONS 0 9731>
 "00000000000000000010011000000100", -- 9731 FREE #<CONS 0 9732>
 "00000000000000000010011000000101", -- 9732 FREE #<CONS 0 9733>
 "00000000000000000010011000000110", -- 9733 FREE #<CONS 0 9734>
 "00000000000000000010011000000111", -- 9734 FREE #<CONS 0 9735>
 "00000000000000000010011000001000", -- 9735 FREE #<CONS 0 9736>
 "00000000000000000010011000001001", -- 9736 FREE #<CONS 0 9737>
 "00000000000000000010011000001010", -- 9737 FREE #<CONS 0 9738>
 "00000000000000000010011000001011", -- 9738 FREE #<CONS 0 9739>
 "00000000000000000010011000001100", -- 9739 FREE #<CONS 0 9740>
 "00000000000000000010011000001101", -- 9740 FREE #<CONS 0 9741>
 "00000000000000000010011000001110", -- 9741 FREE #<CONS 0 9742>
 "00000000000000000010011000001111", -- 9742 FREE #<CONS 0 9743>
 "00000000000000000010011000010000", -- 9743 FREE #<CONS 0 9744>
 "00000000000000000010011000010001", -- 9744 FREE #<CONS 0 9745>
 "00000000000000000010011000010010", -- 9745 FREE #<CONS 0 9746>
 "00000000000000000010011000010011", -- 9746 FREE #<CONS 0 9747>
 "00000000000000000010011000010100", -- 9747 FREE #<CONS 0 9748>
 "00000000000000000010011000010101", -- 9748 FREE #<CONS 0 9749>
 "00000000000000000010011000010110", -- 9749 FREE #<CONS 0 9750>
 "00000000000000000010011000010111", -- 9750 FREE #<CONS 0 9751>
 "00000000000000000010011000011000", -- 9751 FREE #<CONS 0 9752>
 "00000000000000000010011000011001", -- 9752 FREE #<CONS 0 9753>
 "00000000000000000010011000011010", -- 9753 FREE #<CONS 0 9754>
 "00000000000000000010011000011011", -- 9754 FREE #<CONS 0 9755>
 "00000000000000000010011000011100", -- 9755 FREE #<CONS 0 9756>
 "00000000000000000010011000011101", -- 9756 FREE #<CONS 0 9757>
 "00000000000000000010011000011110", -- 9757 FREE #<CONS 0 9758>
 "00000000000000000010011000011111", -- 9758 FREE #<CONS 0 9759>
 "00000000000000000010011000100000", -- 9759 FREE #<CONS 0 9760>
 "00000000000000000010011000100001", -- 9760 FREE #<CONS 0 9761>
 "00000000000000000010011000100010", -- 9761 FREE #<CONS 0 9762>
 "00000000000000000010011000100011", -- 9762 FREE #<CONS 0 9763>
 "00000000000000000010011000100100", -- 9763 FREE #<CONS 0 9764>
 "00000000000000000010011000100101", -- 9764 FREE #<CONS 0 9765>
 "00000000000000000010011000100110", -- 9765 FREE #<CONS 0 9766>
 "00000000000000000010011000100111", -- 9766 FREE #<CONS 0 9767>
 "00000000000000000010011000101000", -- 9767 FREE #<CONS 0 9768>
 "00000000000000000010011000101001", -- 9768 FREE #<CONS 0 9769>
 "00000000000000000010011000101010", -- 9769 FREE #<CONS 0 9770>
 "00000000000000000010011000101011", -- 9770 FREE #<CONS 0 9771>
 "00000000000000000010011000101100", -- 9771 FREE #<CONS 0 9772>
 "00000000000000000010011000101101", -- 9772 FREE #<CONS 0 9773>
 "00000000000000000010011000101110", -- 9773 FREE #<CONS 0 9774>
 "00000000000000000010011000101111", -- 9774 FREE #<CONS 0 9775>
 "00000000000000000010011000110000", -- 9775 FREE #<CONS 0 9776>
 "00000000000000000010011000110001", -- 9776 FREE #<CONS 0 9777>
 "00000000000000000010011000110010", -- 9777 FREE #<CONS 0 9778>
 "00000000000000000010011000110011", -- 9778 FREE #<CONS 0 9779>
 "00000000000000000010011000110100", -- 9779 FREE #<CONS 0 9780>
 "00000000000000000010011000110101", -- 9780 FREE #<CONS 0 9781>
 "00000000000000000010011000110110", -- 9781 FREE #<CONS 0 9782>
 "00000000000000000010011000110111", -- 9782 FREE #<CONS 0 9783>
 "00000000000000000010011000111000", -- 9783 FREE #<CONS 0 9784>
 "00000000000000000010011000111001", -- 9784 FREE #<CONS 0 9785>
 "00000000000000000010011000111010", -- 9785 FREE #<CONS 0 9786>
 "00000000000000000010011000111011", -- 9786 FREE #<CONS 0 9787>
 "00000000000000000010011000111100", -- 9787 FREE #<CONS 0 9788>
 "00000000000000000010011000111101", -- 9788 FREE #<CONS 0 9789>
 "00000000000000000010011000111110", -- 9789 FREE #<CONS 0 9790>
 "00000000000000000010011000111111", -- 9790 FREE #<CONS 0 9791>
 "00000000000000000010011001000000", -- 9791 FREE #<CONS 0 9792>
 "00000000000000000010011001000001", -- 9792 FREE #<CONS 0 9793>
 "00000000000000000010011001000010", -- 9793 FREE #<CONS 0 9794>
 "00000000000000000010011001000011", -- 9794 FREE #<CONS 0 9795>
 "00000000000000000010011001000100", -- 9795 FREE #<CONS 0 9796>
 "00000000000000000010011001000101", -- 9796 FREE #<CONS 0 9797>
 "00000000000000000010011001000110", -- 9797 FREE #<CONS 0 9798>
 "00000000000000000010011001000111", -- 9798 FREE #<CONS 0 9799>
 "00000000000000000010011001001000", -- 9799 FREE #<CONS 0 9800>
 "00000000000000000010011001001001", -- 9800 FREE #<CONS 0 9801>
 "00000000000000000010011001001010", -- 9801 FREE #<CONS 0 9802>
 "00000000000000000010011001001011", -- 9802 FREE #<CONS 0 9803>
 "00000000000000000010011001001100", -- 9803 FREE #<CONS 0 9804>
 "00000000000000000010011001001101", -- 9804 FREE #<CONS 0 9805>
 "00000000000000000010011001001110", -- 9805 FREE #<CONS 0 9806>
 "00000000000000000010011001001111", -- 9806 FREE #<CONS 0 9807>
 "00000000000000000010011001010000", -- 9807 FREE #<CONS 0 9808>
 "00000000000000000010011001010001", -- 9808 FREE #<CONS 0 9809>
 "00000000000000000010011001010010", -- 9809 FREE #<CONS 0 9810>
 "00000000000000000010011001010011", -- 9810 FREE #<CONS 0 9811>
 "00000000000000000010011001010100", -- 9811 FREE #<CONS 0 9812>
 "00000000000000000010011001010101", -- 9812 FREE #<CONS 0 9813>
 "00000000000000000010011001010110", -- 9813 FREE #<CONS 0 9814>
 "00000000000000000010011001010111", -- 9814 FREE #<CONS 0 9815>
 "00000000000000000010011001011000", -- 9815 FREE #<CONS 0 9816>
 "00000000000000000010011001011001", -- 9816 FREE #<CONS 0 9817>
 "00000000000000000010011001011010", -- 9817 FREE #<CONS 0 9818>
 "00000000000000000010011001011011", -- 9818 FREE #<CONS 0 9819>
 "00000000000000000010011001011100", -- 9819 FREE #<CONS 0 9820>
 "00000000000000000010011001011101", -- 9820 FREE #<CONS 0 9821>
 "00000000000000000010011001011110", -- 9821 FREE #<CONS 0 9822>
 "00000000000000000010011001011111", -- 9822 FREE #<CONS 0 9823>
 "00000000000000000010011001100000", -- 9823 FREE #<CONS 0 9824>
 "00000000000000000010011001100001", -- 9824 FREE #<CONS 0 9825>
 "00000000000000000010011001100010", -- 9825 FREE #<CONS 0 9826>
 "00000000000000000010011001100011", -- 9826 FREE #<CONS 0 9827>
 "00000000000000000010011001100100", -- 9827 FREE #<CONS 0 9828>
 "00000000000000000010011001100101", -- 9828 FREE #<CONS 0 9829>
 "00000000000000000010011001100110", -- 9829 FREE #<CONS 0 9830>
 "00000000000000000010011001100111", -- 9830 FREE #<CONS 0 9831>
 "00000000000000000010011001101000", -- 9831 FREE #<CONS 0 9832>
 "00000000000000000010011001101001", -- 9832 FREE #<CONS 0 9833>
 "00000000000000000010011001101010", -- 9833 FREE #<CONS 0 9834>
 "00000000000000000010011001101011", -- 9834 FREE #<CONS 0 9835>
 "00000000000000000010011001101100", -- 9835 FREE #<CONS 0 9836>
 "00000000000000000010011001101101", -- 9836 FREE #<CONS 0 9837>
 "00000000000000000010011001101110", -- 9837 FREE #<CONS 0 9838>
 "00000000000000000010011001101111", -- 9838 FREE #<CONS 0 9839>
 "00000000000000000010011001110000", -- 9839 FREE #<CONS 0 9840>
 "00000000000000000010011001110001", -- 9840 FREE #<CONS 0 9841>
 "00000000000000000010011001110010", -- 9841 FREE #<CONS 0 9842>
 "00000000000000000010011001110011", -- 9842 FREE #<CONS 0 9843>
 "00000000000000000010011001110100", -- 9843 FREE #<CONS 0 9844>
 "00000000000000000010011001110101", -- 9844 FREE #<CONS 0 9845>
 "00000000000000000010011001110110", -- 9845 FREE #<CONS 0 9846>
 "00000000000000000010011001110111", -- 9846 FREE #<CONS 0 9847>
 "00000000000000000010011001111000", -- 9847 FREE #<CONS 0 9848>
 "00000000000000000010011001111001", -- 9848 FREE #<CONS 0 9849>
 "00000000000000000010011001111010", -- 9849 FREE #<CONS 0 9850>
 "00000000000000000010011001111011", -- 9850 FREE #<CONS 0 9851>
 "00000000000000000010011001111100", -- 9851 FREE #<CONS 0 9852>
 "00000000000000000010011001111101", -- 9852 FREE #<CONS 0 9853>
 "00000000000000000010011001111110", -- 9853 FREE #<CONS 0 9854>
 "00000000000000000010011001111111", -- 9854 FREE #<CONS 0 9855>
 "00000000000000000010011010000000", -- 9855 FREE #<CONS 0 9856>
 "00000000000000000010011010000001", -- 9856 FREE #<CONS 0 9857>
 "00000000000000000010011010000010", -- 9857 FREE #<CONS 0 9858>
 "00000000000000000010011010000011", -- 9858 FREE #<CONS 0 9859>
 "00000000000000000010011010000100", -- 9859 FREE #<CONS 0 9860>
 "00000000000000000010011010000101", -- 9860 FREE #<CONS 0 9861>
 "00000000000000000010011010000110", -- 9861 FREE #<CONS 0 9862>
 "00000000000000000010011010000111", -- 9862 FREE #<CONS 0 9863>
 "00000000000000000010011010001000", -- 9863 FREE #<CONS 0 9864>
 "00000000000000000010011010001001", -- 9864 FREE #<CONS 0 9865>
 "00000000000000000010011010001010", -- 9865 FREE #<CONS 0 9866>
 "00000000000000000010011010001011", -- 9866 FREE #<CONS 0 9867>
 "00000000000000000010011010001100", -- 9867 FREE #<CONS 0 9868>
 "00000000000000000010011010001101", -- 9868 FREE #<CONS 0 9869>
 "00000000000000000010011010001110", -- 9869 FREE #<CONS 0 9870>
 "00000000000000000010011010001111", -- 9870 FREE #<CONS 0 9871>
 "00000000000000000010011010010000", -- 9871 FREE #<CONS 0 9872>
 "00000000000000000010011010010001", -- 9872 FREE #<CONS 0 9873>
 "00000000000000000010011010010010", -- 9873 FREE #<CONS 0 9874>
 "00000000000000000010011010010011", -- 9874 FREE #<CONS 0 9875>
 "00000000000000000010011010010100", -- 9875 FREE #<CONS 0 9876>
 "00000000000000000010011010010101", -- 9876 FREE #<CONS 0 9877>
 "00000000000000000010011010010110", -- 9877 FREE #<CONS 0 9878>
 "00000000000000000010011010010111", -- 9878 FREE #<CONS 0 9879>
 "00000000000000000010011010011000", -- 9879 FREE #<CONS 0 9880>
 "00000000000000000010011010011001", -- 9880 FREE #<CONS 0 9881>
 "00000000000000000010011010011010", -- 9881 FREE #<CONS 0 9882>
 "00000000000000000010011010011011", -- 9882 FREE #<CONS 0 9883>
 "00000000000000000010011010011100", -- 9883 FREE #<CONS 0 9884>
 "00000000000000000010011010011101", -- 9884 FREE #<CONS 0 9885>
 "00000000000000000010011010011110", -- 9885 FREE #<CONS 0 9886>
 "00000000000000000010011010011111", -- 9886 FREE #<CONS 0 9887>
 "00000000000000000010011010100000", -- 9887 FREE #<CONS 0 9888>
 "00000000000000000010011010100001", -- 9888 FREE #<CONS 0 9889>
 "00000000000000000010011010100010", -- 9889 FREE #<CONS 0 9890>
 "00000000000000000010011010100011", -- 9890 FREE #<CONS 0 9891>
 "00000000000000000010011010100100", -- 9891 FREE #<CONS 0 9892>
 "00000000000000000010011010100101", -- 9892 FREE #<CONS 0 9893>
 "00000000000000000010011010100110", -- 9893 FREE #<CONS 0 9894>
 "00000000000000000010011010100111", -- 9894 FREE #<CONS 0 9895>
 "00000000000000000010011010101000", -- 9895 FREE #<CONS 0 9896>
 "00000000000000000010011010101001", -- 9896 FREE #<CONS 0 9897>
 "00000000000000000010011010101010", -- 9897 FREE #<CONS 0 9898>
 "00000000000000000010011010101011", -- 9898 FREE #<CONS 0 9899>
 "00000000000000000010011010101100", -- 9899 FREE #<CONS 0 9900>
 "00000000000000000010011010101101", -- 9900 FREE #<CONS 0 9901>
 "00000000000000000010011010101110", -- 9901 FREE #<CONS 0 9902>
 "00000000000000000010011010101111", -- 9902 FREE #<CONS 0 9903>
 "00000000000000000010011010110000", -- 9903 FREE #<CONS 0 9904>
 "00000000000000000010011010110001", -- 9904 FREE #<CONS 0 9905>
 "00000000000000000010011010110010", -- 9905 FREE #<CONS 0 9906>
 "00000000000000000010011010110011", -- 9906 FREE #<CONS 0 9907>
 "00000000000000000010011010110100", -- 9907 FREE #<CONS 0 9908>
 "00000000000000000010011010110101", -- 9908 FREE #<CONS 0 9909>
 "00000000000000000010011010110110", -- 9909 FREE #<CONS 0 9910>
 "00000000000000000010011010110111", -- 9910 FREE #<CONS 0 9911>
 "00000000000000000010011010111000", -- 9911 FREE #<CONS 0 9912>
 "00000000000000000010011010111001", -- 9912 FREE #<CONS 0 9913>
 "00000000000000000010011010111010", -- 9913 FREE #<CONS 0 9914>
 "00000000000000000010011010111011", -- 9914 FREE #<CONS 0 9915>
 "00000000000000000010011010111100", -- 9915 FREE #<CONS 0 9916>
 "00000000000000000010011010111101", -- 9916 FREE #<CONS 0 9917>
 "00000000000000000010011010111110", -- 9917 FREE #<CONS 0 9918>
 "00000000000000000010011010111111", -- 9918 FREE #<CONS 0 9919>
 "00000000000000000010011011000000", -- 9919 FREE #<CONS 0 9920>
 "00000000000000000010011011000001", -- 9920 FREE #<CONS 0 9921>
 "00000000000000000010011011000010", -- 9921 FREE #<CONS 0 9922>
 "00000000000000000010011011000011", -- 9922 FREE #<CONS 0 9923>
 "00000000000000000010011011000100", -- 9923 FREE #<CONS 0 9924>
 "00000000000000000010011011000101", -- 9924 FREE #<CONS 0 9925>
 "00000000000000000010011011000110", -- 9925 FREE #<CONS 0 9926>
 "00000000000000000010011011000111", -- 9926 FREE #<CONS 0 9927>
 "00000000000000000010011011001000", -- 9927 FREE #<CONS 0 9928>
 "00000000000000000010011011001001", -- 9928 FREE #<CONS 0 9929>
 "00000000000000000010011011001010", -- 9929 FREE #<CONS 0 9930>
 "00000000000000000010011011001011", -- 9930 FREE #<CONS 0 9931>
 "00000000000000000010011011001100", -- 9931 FREE #<CONS 0 9932>
 "00000000000000000010011011001101", -- 9932 FREE #<CONS 0 9933>
 "00000000000000000010011011001110", -- 9933 FREE #<CONS 0 9934>
 "00000000000000000010011011001111", -- 9934 FREE #<CONS 0 9935>
 "00000000000000000010011011010000", -- 9935 FREE #<CONS 0 9936>
 "00000000000000000010011011010001", -- 9936 FREE #<CONS 0 9937>
 "00000000000000000010011011010010", -- 9937 FREE #<CONS 0 9938>
 "00000000000000000010011011010011", -- 9938 FREE #<CONS 0 9939>
 "00000000000000000010011011010100", -- 9939 FREE #<CONS 0 9940>
 "00000000000000000010011011010101", -- 9940 FREE #<CONS 0 9941>
 "00000000000000000010011011010110", -- 9941 FREE #<CONS 0 9942>
 "00000000000000000010011011010111", -- 9942 FREE #<CONS 0 9943>
 "00000000000000000010011011011000", -- 9943 FREE #<CONS 0 9944>
 "00000000000000000010011011011001", -- 9944 FREE #<CONS 0 9945>
 "00000000000000000010011011011010", -- 9945 FREE #<CONS 0 9946>
 "00000000000000000010011011011011", -- 9946 FREE #<CONS 0 9947>
 "00000000000000000010011011011100", -- 9947 FREE #<CONS 0 9948>
 "00000000000000000010011011011101", -- 9948 FREE #<CONS 0 9949>
 "00000000000000000010011011011110", -- 9949 FREE #<CONS 0 9950>
 "00000000000000000010011011011111", -- 9950 FREE #<CONS 0 9951>
 "00000000000000000010011011100000", -- 9951 FREE #<CONS 0 9952>
 "00000000000000000010011011100001", -- 9952 FREE #<CONS 0 9953>
 "00000000000000000010011011100010", -- 9953 FREE #<CONS 0 9954>
 "00000000000000000010011011100011", -- 9954 FREE #<CONS 0 9955>
 "00000000000000000010011011100100", -- 9955 FREE #<CONS 0 9956>
 "00000000000000000010011011100101", -- 9956 FREE #<CONS 0 9957>
 "00000000000000000010011011100110", -- 9957 FREE #<CONS 0 9958>
 "00000000000000000010011011100111", -- 9958 FREE #<CONS 0 9959>
 "00000000000000000010011011101000", -- 9959 FREE #<CONS 0 9960>
 "00000000000000000010011011101001", -- 9960 FREE #<CONS 0 9961>
 "00000000000000000010011011101010", -- 9961 FREE #<CONS 0 9962>
 "00000000000000000010011011101011", -- 9962 FREE #<CONS 0 9963>
 "00000000000000000010011011101100", -- 9963 FREE #<CONS 0 9964>
 "00000000000000000010011011101101", -- 9964 FREE #<CONS 0 9965>
 "00000000000000000010011011101110", -- 9965 FREE #<CONS 0 9966>
 "00000000000000000010011011101111", -- 9966 FREE #<CONS 0 9967>
 "00000000000000000010011011110000", -- 9967 FREE #<CONS 0 9968>
 "00000000000000000010011011110001", -- 9968 FREE #<CONS 0 9969>
 "00000000000000000010011011110010", -- 9969 FREE #<CONS 0 9970>
 "00000000000000000010011011110011", -- 9970 FREE #<CONS 0 9971>
 "00000000000000000010011011110100", -- 9971 FREE #<CONS 0 9972>
 "00000000000000000010011011110101", -- 9972 FREE #<CONS 0 9973>
 "00000000000000000010011011110110", -- 9973 FREE #<CONS 0 9974>
 "00000000000000000010011011110111", -- 9974 FREE #<CONS 0 9975>
 "00000000000000000010011011111000", -- 9975 FREE #<CONS 0 9976>
 "00000000000000000010011011111001", -- 9976 FREE #<CONS 0 9977>
 "00000000000000000010011011111010", -- 9977 FREE #<CONS 0 9978>
 "00000000000000000010011011111011", -- 9978 FREE #<CONS 0 9979>
 "00000000000000000010011011111100", -- 9979 FREE #<CONS 0 9980>
 "00000000000000000010011011111101", -- 9980 FREE #<CONS 0 9981>
 "00000000000000000010011011111110", -- 9981 FREE #<CONS 0 9982>
 "00000000000000000010011011111111", -- 9982 FREE #<CONS 0 9983>
 "00000000000000000010011100000000", -- 9983 FREE #<CONS 0 9984>
 "00000000000000000010011100000001", -- 9984 FREE #<CONS 0 9985>
 "00000000000000000010011100000010", -- 9985 FREE #<CONS 0 9986>
 "00000000000000000010011100000011", -- 9986 FREE #<CONS 0 9987>
 "00000000000000000010011100000100", -- 9987 FREE #<CONS 0 9988>
 "00000000000000000010011100000101", -- 9988 FREE #<CONS 0 9989>
 "00000000000000000010011100000110", -- 9989 FREE #<CONS 0 9990>
 "00000000000000000010011100000111", -- 9990 FREE #<CONS 0 9991>
 "00000000000000000010011100001000", -- 9991 FREE #<CONS 0 9992>
 "00000000000000000010011100001001", -- 9992 FREE #<CONS 0 9993>
 "00000000000000000010011100001010", -- 9993 FREE #<CONS 0 9994>
 "00000000000000000010011100001011", -- 9994 FREE #<CONS 0 9995>
 "00000000000000000010011100001100", -- 9995 FREE #<CONS 0 9996>
 "00000000000000000010011100001101", -- 9996 FREE #<CONS 0 9997>
 "00000000000000000010011100001110", -- 9997 FREE #<CONS 0 9998>
 "00000000000000000010011100001111", -- 9998 FREE #<CONS 0 9999>
 "00000000000000000010011100010000", -- 9999 FREE #<CONS 0 10000>
 "00000000000000000010011100010001", -- 10000 FREE #<CONS 0 10001>
 "00000000000000000010011100010010", -- 10001 FREE #<CONS 0 10002>
 "00000000000000000010011100010011", -- 10002 FREE #<CONS 0 10003>
 "00000000000000000010011100010100", -- 10003 FREE #<CONS 0 10004>
 "00000000000000000010011100010101", -- 10004 FREE #<CONS 0 10005>
 "00000000000000000010011100010110", -- 10005 FREE #<CONS 0 10006>
 "00000000000000000010011100010111", -- 10006 FREE #<CONS 0 10007>
 "00000000000000000010011100011000", -- 10007 FREE #<CONS 0 10008>
 "00000000000000000010011100011001", -- 10008 FREE #<CONS 0 10009>
 "00000000000000000010011100011010", -- 10009 FREE #<CONS 0 10010>
 "00000000000000000010011100011011", -- 10010 FREE #<CONS 0 10011>
 "00000000000000000010011100011100", -- 10011 FREE #<CONS 0 10012>
 "00000000000000000010011100011101", -- 10012 FREE #<CONS 0 10013>
 "00000000000000000010011100011110", -- 10013 FREE #<CONS 0 10014>
 "00000000000000000010011100011111", -- 10014 FREE #<CONS 0 10015>
 "00000000000000000010011100100000", -- 10015 FREE #<CONS 0 10016>
 "00000000000000000010011100100001", -- 10016 FREE #<CONS 0 10017>
 "00000000000000000010011100100010", -- 10017 FREE #<CONS 0 10018>
 "00000000000000000010011100100011", -- 10018 FREE #<CONS 0 10019>
 "00000000000000000010011100100100", -- 10019 FREE #<CONS 0 10020>
 "00000000000000000010011100100101", -- 10020 FREE #<CONS 0 10021>
 "00000000000000000010011100100110", -- 10021 FREE #<CONS 0 10022>
 "00000000000000000010011100100111", -- 10022 FREE #<CONS 0 10023>
 "00000000000000000010011100101000", -- 10023 FREE #<CONS 0 10024>
 "00000000000000000010011100101001", -- 10024 FREE #<CONS 0 10025>
 "00000000000000000010011100101010", -- 10025 FREE #<CONS 0 10026>
 "00000000000000000010011100101011", -- 10026 FREE #<CONS 0 10027>
 "00000000000000000010011100101100", -- 10027 FREE #<CONS 0 10028>
 "00000000000000000010011100101101", -- 10028 FREE #<CONS 0 10029>
 "00000000000000000010011100101110", -- 10029 FREE #<CONS 0 10030>
 "00000000000000000010011100101111", -- 10030 FREE #<CONS 0 10031>
 "00000000000000000010011100110000", -- 10031 FREE #<CONS 0 10032>
 "00000000000000000010011100110001", -- 10032 FREE #<CONS 0 10033>
 "00000000000000000010011100110010", -- 10033 FREE #<CONS 0 10034>
 "00000000000000000010011100110011", -- 10034 FREE #<CONS 0 10035>
 "00000000000000000010011100110100", -- 10035 FREE #<CONS 0 10036>
 "00000000000000000010011100110101", -- 10036 FREE #<CONS 0 10037>
 "00000000000000000010011100110110", -- 10037 FREE #<CONS 0 10038>
 "00000000000000000010011100110111", -- 10038 FREE #<CONS 0 10039>
 "00000000000000000010011100111000", -- 10039 FREE #<CONS 0 10040>
 "00000000000000000010011100111001", -- 10040 FREE #<CONS 0 10041>
 "00000000000000000010011100111010", -- 10041 FREE #<CONS 0 10042>
 "00000000000000000010011100111011", -- 10042 FREE #<CONS 0 10043>
 "00000000000000000010011100111100", -- 10043 FREE #<CONS 0 10044>
 "00000000000000000010011100111101", -- 10044 FREE #<CONS 0 10045>
 "00000000000000000010011100111110", -- 10045 FREE #<CONS 0 10046>
 "00000000000000000010011100111111", -- 10046 FREE #<CONS 0 10047>
 "00000000000000000010011101000000", -- 10047 FREE #<CONS 0 10048>
 "00000000000000000010011101000001", -- 10048 FREE #<CONS 0 10049>
 "00000000000000000010011101000010", -- 10049 FREE #<CONS 0 10050>
 "00000000000000000010011101000011", -- 10050 FREE #<CONS 0 10051>
 "00000000000000000010011101000100", -- 10051 FREE #<CONS 0 10052>
 "00000000000000000010011101000101", -- 10052 FREE #<CONS 0 10053>
 "00000000000000000010011101000110", -- 10053 FREE #<CONS 0 10054>
 "00000000000000000010011101000111", -- 10054 FREE #<CONS 0 10055>
 "00000000000000000010011101001000", -- 10055 FREE #<CONS 0 10056>
 "00000000000000000010011101001001", -- 10056 FREE #<CONS 0 10057>
 "00000000000000000010011101001010", -- 10057 FREE #<CONS 0 10058>
 "00000000000000000010011101001011", -- 10058 FREE #<CONS 0 10059>
 "00000000000000000010011101001100", -- 10059 FREE #<CONS 0 10060>
 "00000000000000000010011101001101", -- 10060 FREE #<CONS 0 10061>
 "00000000000000000010011101001110", -- 10061 FREE #<CONS 0 10062>
 "00000000000000000010011101001111", -- 10062 FREE #<CONS 0 10063>
 "00000000000000000010011101010000", -- 10063 FREE #<CONS 0 10064>
 "00000000000000000010011101010001", -- 10064 FREE #<CONS 0 10065>
 "00000000000000000010011101010010", -- 10065 FREE #<CONS 0 10066>
 "00000000000000000010011101010011", -- 10066 FREE #<CONS 0 10067>
 "00000000000000000010011101010100", -- 10067 FREE #<CONS 0 10068>
 "00000000000000000010011101010101", -- 10068 FREE #<CONS 0 10069>
 "00000000000000000010011101010110", -- 10069 FREE #<CONS 0 10070>
 "00000000000000000010011101010111", -- 10070 FREE #<CONS 0 10071>
 "00000000000000000010011101011000", -- 10071 FREE #<CONS 0 10072>
 "00000000000000000010011101011001", -- 10072 FREE #<CONS 0 10073>
 "00000000000000000010011101011010", -- 10073 FREE #<CONS 0 10074>
 "00000000000000000010011101011011", -- 10074 FREE #<CONS 0 10075>
 "00000000000000000010011101011100", -- 10075 FREE #<CONS 0 10076>
 "00000000000000000010011101011101", -- 10076 FREE #<CONS 0 10077>
 "00000000000000000010011101011110", -- 10077 FREE #<CONS 0 10078>
 "00000000000000000010011101011111", -- 10078 FREE #<CONS 0 10079>
 "00000000000000000010011101100000", -- 10079 FREE #<CONS 0 10080>
 "00000000000000000010011101100001", -- 10080 FREE #<CONS 0 10081>
 "00000000000000000010011101100010", -- 10081 FREE #<CONS 0 10082>
 "00000000000000000010011101100011", -- 10082 FREE #<CONS 0 10083>
 "00000000000000000010011101100100", -- 10083 FREE #<CONS 0 10084>
 "00000000000000000010011101100101", -- 10084 FREE #<CONS 0 10085>
 "00000000000000000010011101100110", -- 10085 FREE #<CONS 0 10086>
 "00000000000000000010011101100111", -- 10086 FREE #<CONS 0 10087>
 "00000000000000000010011101101000", -- 10087 FREE #<CONS 0 10088>
 "00000000000000000010011101101001", -- 10088 FREE #<CONS 0 10089>
 "00000000000000000010011101101010", -- 10089 FREE #<CONS 0 10090>
 "00000000000000000010011101101011", -- 10090 FREE #<CONS 0 10091>
 "00000000000000000010011101101100", -- 10091 FREE #<CONS 0 10092>
 "00000000000000000010011101101101", -- 10092 FREE #<CONS 0 10093>
 "00000000000000000010011101101110", -- 10093 FREE #<CONS 0 10094>
 "00000000000000000010011101101111", -- 10094 FREE #<CONS 0 10095>
 "00000000000000000010011101110000", -- 10095 FREE #<CONS 0 10096>
 "00000000000000000010011101110001", -- 10096 FREE #<CONS 0 10097>
 "00000000000000000010011101110010", -- 10097 FREE #<CONS 0 10098>
 "00000000000000000010011101110011", -- 10098 FREE #<CONS 0 10099>
 "00000000000000000010011101110100", -- 10099 FREE #<CONS 0 10100>
 "00000000000000000010011101110101", -- 10100 FREE #<CONS 0 10101>
 "00000000000000000010011101110110", -- 10101 FREE #<CONS 0 10102>
 "00000000000000000010011101110111", -- 10102 FREE #<CONS 0 10103>
 "00000000000000000010011101111000", -- 10103 FREE #<CONS 0 10104>
 "00000000000000000010011101111001", -- 10104 FREE #<CONS 0 10105>
 "00000000000000000010011101111010", -- 10105 FREE #<CONS 0 10106>
 "00000000000000000010011101111011", -- 10106 FREE #<CONS 0 10107>
 "00000000000000000010011101111100", -- 10107 FREE #<CONS 0 10108>
 "00000000000000000010011101111101", -- 10108 FREE #<CONS 0 10109>
 "00000000000000000010011101111110", -- 10109 FREE #<CONS 0 10110>
 "00000000000000000010011101111111", -- 10110 FREE #<CONS 0 10111>
 "00000000000000000010011110000000", -- 10111 FREE #<CONS 0 10112>
 "00000000000000000010011110000001", -- 10112 FREE #<CONS 0 10113>
 "00000000000000000010011110000010", -- 10113 FREE #<CONS 0 10114>
 "00000000000000000010011110000011", -- 10114 FREE #<CONS 0 10115>
 "00000000000000000010011110000100", -- 10115 FREE #<CONS 0 10116>
 "00000000000000000010011110000101", -- 10116 FREE #<CONS 0 10117>
 "00000000000000000010011110000110", -- 10117 FREE #<CONS 0 10118>
 "00000000000000000010011110000111", -- 10118 FREE #<CONS 0 10119>
 "00000000000000000010011110001000", -- 10119 FREE #<CONS 0 10120>
 "00000000000000000010011110001001", -- 10120 FREE #<CONS 0 10121>
 "00000000000000000010011110001010", -- 10121 FREE #<CONS 0 10122>
 "00000000000000000010011110001011", -- 10122 FREE #<CONS 0 10123>
 "00000000000000000010011110001100", -- 10123 FREE #<CONS 0 10124>
 "00000000000000000010011110001101", -- 10124 FREE #<CONS 0 10125>
 "00000000000000000010011110001110", -- 10125 FREE #<CONS 0 10126>
 "00000000000000000010011110001111", -- 10126 FREE #<CONS 0 10127>
 "00000000000000000010011110010000", -- 10127 FREE #<CONS 0 10128>
 "00000000000000000010011110010001", -- 10128 FREE #<CONS 0 10129>
 "00000000000000000010011110010010", -- 10129 FREE #<CONS 0 10130>
 "00000000000000000010011110010011", -- 10130 FREE #<CONS 0 10131>
 "00000000000000000010011110010100", -- 10131 FREE #<CONS 0 10132>
 "00000000000000000010011110010101", -- 10132 FREE #<CONS 0 10133>
 "00000000000000000010011110010110", -- 10133 FREE #<CONS 0 10134>
 "00000000000000000010011110010111", -- 10134 FREE #<CONS 0 10135>
 "00000000000000000010011110011000", -- 10135 FREE #<CONS 0 10136>
 "00000000000000000010011110011001", -- 10136 FREE #<CONS 0 10137>
 "00000000000000000010011110011010", -- 10137 FREE #<CONS 0 10138>
 "00000000000000000010011110011011", -- 10138 FREE #<CONS 0 10139>
 "00000000000000000010011110011100", -- 10139 FREE #<CONS 0 10140>
 "00000000000000000010011110011101", -- 10140 FREE #<CONS 0 10141>
 "00000000000000000010011110011110", -- 10141 FREE #<CONS 0 10142>
 "00000000000000000010011110011111", -- 10142 FREE #<CONS 0 10143>
 "00000000000000000010011110100000", -- 10143 FREE #<CONS 0 10144>
 "00000000000000000010011110100001", -- 10144 FREE #<CONS 0 10145>
 "00000000000000000010011110100010", -- 10145 FREE #<CONS 0 10146>
 "00000000000000000010011110100011", -- 10146 FREE #<CONS 0 10147>
 "00000000000000000010011110100100", -- 10147 FREE #<CONS 0 10148>
 "00000000000000000010011110100101", -- 10148 FREE #<CONS 0 10149>
 "00000000000000000010011110100110", -- 10149 FREE #<CONS 0 10150>
 "00000000000000000010011110100111", -- 10150 FREE #<CONS 0 10151>
 "00000000000000000010011110101000", -- 10151 FREE #<CONS 0 10152>
 "00000000000000000010011110101001", -- 10152 FREE #<CONS 0 10153>
 "00000000000000000010011110101010", -- 10153 FREE #<CONS 0 10154>
 "00000000000000000010011110101011", -- 10154 FREE #<CONS 0 10155>
 "00000000000000000010011110101100", -- 10155 FREE #<CONS 0 10156>
 "00000000000000000010011110101101", -- 10156 FREE #<CONS 0 10157>
 "00000000000000000010011110101110", -- 10157 FREE #<CONS 0 10158>
 "00000000000000000010011110101111", -- 10158 FREE #<CONS 0 10159>
 "00000000000000000010011110110000", -- 10159 FREE #<CONS 0 10160>
 "00000000000000000010011110110001", -- 10160 FREE #<CONS 0 10161>
 "00000000000000000010011110110010", -- 10161 FREE #<CONS 0 10162>
 "00000000000000000010011110110011", -- 10162 FREE #<CONS 0 10163>
 "00000000000000000010011110110100", -- 10163 FREE #<CONS 0 10164>
 "00000000000000000010011110110101", -- 10164 FREE #<CONS 0 10165>
 "00000000000000000010011110110110", -- 10165 FREE #<CONS 0 10166>
 "00000000000000000010011110110111", -- 10166 FREE #<CONS 0 10167>
 "00000000000000000010011110111000", -- 10167 FREE #<CONS 0 10168>
 "00000000000000000010011110111001", -- 10168 FREE #<CONS 0 10169>
 "00000000000000000010011110111010", -- 10169 FREE #<CONS 0 10170>
 "00000000000000000010011110111011", -- 10170 FREE #<CONS 0 10171>
 "00000000000000000010011110111100", -- 10171 FREE #<CONS 0 10172>
 "00000000000000000010011110111101", -- 10172 FREE #<CONS 0 10173>
 "00000000000000000010011110111110", -- 10173 FREE #<CONS 0 10174>
 "00000000000000000010011110111111", -- 10174 FREE #<CONS 0 10175>
 "00000000000000000010011111000000", -- 10175 FREE #<CONS 0 10176>
 "00000000000000000010011111000001", -- 10176 FREE #<CONS 0 10177>
 "00000000000000000010011111000010", -- 10177 FREE #<CONS 0 10178>
 "00000000000000000010011111000011", -- 10178 FREE #<CONS 0 10179>
 "00000000000000000010011111000100", -- 10179 FREE #<CONS 0 10180>
 "00000000000000000010011111000101", -- 10180 FREE #<CONS 0 10181>
 "00000000000000000010011111000110", -- 10181 FREE #<CONS 0 10182>
 "00000000000000000010011111000111", -- 10182 FREE #<CONS 0 10183>
 "00000000000000000010011111001000", -- 10183 FREE #<CONS 0 10184>
 "00000000000000000010011111001001", -- 10184 FREE #<CONS 0 10185>
 "00000000000000000010011111001010", -- 10185 FREE #<CONS 0 10186>
 "00000000000000000010011111001011", -- 10186 FREE #<CONS 0 10187>
 "00000000000000000010011111001100", -- 10187 FREE #<CONS 0 10188>
 "00000000000000000010011111001101", -- 10188 FREE #<CONS 0 10189>
 "00000000000000000010011111001110", -- 10189 FREE #<CONS 0 10190>
 "00000000000000000010011111001111", -- 10190 FREE #<CONS 0 10191>
 "00000000000000000010011111010000", -- 10191 FREE #<CONS 0 10192>
 "00000000000000000010011111010001", -- 10192 FREE #<CONS 0 10193>
 "00000000000000000010011111010010", -- 10193 FREE #<CONS 0 10194>
 "00000000000000000010011111010011", -- 10194 FREE #<CONS 0 10195>
 "00000000000000000010011111010100", -- 10195 FREE #<CONS 0 10196>
 "00000000000000000010011111010101", -- 10196 FREE #<CONS 0 10197>
 "00000000000000000010011111010110", -- 10197 FREE #<CONS 0 10198>
 "00000000000000000010011111010111", -- 10198 FREE #<CONS 0 10199>
 "00000000000000000010011111011000", -- 10199 FREE #<CONS 0 10200>
 "00000000000000000010011111011001", -- 10200 FREE #<CONS 0 10201>
 "00000000000000000010011111011010", -- 10201 FREE #<CONS 0 10202>
 "00000000000000000010011111011011", -- 10202 FREE #<CONS 0 10203>
 "00000000000000000010011111011100", -- 10203 FREE #<CONS 0 10204>
 "00000000000000000010011111011101", -- 10204 FREE #<CONS 0 10205>
 "00000000000000000010011111011110", -- 10205 FREE #<CONS 0 10206>
 "00000000000000000010011111011111", -- 10206 FREE #<CONS 0 10207>
 "00000000000000000010011111100000", -- 10207 FREE #<CONS 0 10208>
 "00000000000000000010011111100001", -- 10208 FREE #<CONS 0 10209>
 "00000000000000000010011111100010", -- 10209 FREE #<CONS 0 10210>
 "00000000000000000010011111100011", -- 10210 FREE #<CONS 0 10211>
 "00000000000000000010011111100100", -- 10211 FREE #<CONS 0 10212>
 "00000000000000000010011111100101", -- 10212 FREE #<CONS 0 10213>
 "00000000000000000010011111100110", -- 10213 FREE #<CONS 0 10214>
 "00000000000000000010011111100111", -- 10214 FREE #<CONS 0 10215>
 "00000000000000000010011111101000", -- 10215 FREE #<CONS 0 10216>
 "00000000000000000010011111101001", -- 10216 FREE #<CONS 0 10217>
 "00000000000000000010011111101010", -- 10217 FREE #<CONS 0 10218>
 "00000000000000000010011111101011", -- 10218 FREE #<CONS 0 10219>
 "00000000000000000010011111101100", -- 10219 FREE #<CONS 0 10220>
 "00000000000000000010011111101101", -- 10220 FREE #<CONS 0 10221>
 "00000000000000000010011111101110", -- 10221 FREE #<CONS 0 10222>
 "00000000000000000010011111101111", -- 10222 FREE #<CONS 0 10223>
 "00000000000000000010011111110000", -- 10223 FREE #<CONS 0 10224>
 "00000000000000000010011111110001", -- 10224 FREE #<CONS 0 10225>
 "00000000000000000010011111110010", -- 10225 FREE #<CONS 0 10226>
 "00000000000000000010011111110011", -- 10226 FREE #<CONS 0 10227>
 "00000000000000000010011111110100", -- 10227 FREE #<CONS 0 10228>
 "00000000000000000010011111110101", -- 10228 FREE #<CONS 0 10229>
 "00000000000000000010011111110110", -- 10229 FREE #<CONS 0 10230>
 "00000000000000000010011111110111", -- 10230 FREE #<CONS 0 10231>
 "00000000000000000010011111111000", -- 10231 FREE #<CONS 0 10232>
 "00000000000000000010011111111001", -- 10232 FREE #<CONS 0 10233>
 "00000000000000000010011111111010", -- 10233 FREE #<CONS 0 10234>
 "00000000000000000010011111111011", -- 10234 FREE #<CONS 0 10235>
 "00000000000000000010011111111100", -- 10235 FREE #<CONS 0 10236>
 "00000000000000000010011111111101", -- 10236 FREE #<CONS 0 10237>
 "00000000000000000010011111111110", -- 10237 FREE #<CONS 0 10238>
 "00000000000000000010011111111111", -- 10238 FREE #<CONS 0 10239>
 "00000000000000000010100000000000", -- 10239 FREE #<CONS 0 10240>
 "00000000000000000010100000000001", -- 10240 FREE #<CONS 0 10241>
 "00000000000000000010100000000010", -- 10241 FREE #<CONS 0 10242>
 "00000000000000000010100000000011", -- 10242 FREE #<CONS 0 10243>
 "00000000000000000010100000000100", -- 10243 FREE #<CONS 0 10244>
 "00000000000000000010100000000101", -- 10244 FREE #<CONS 0 10245>
 "00000000000000000010100000000110", -- 10245 FREE #<CONS 0 10246>
 "00000000000000000010100000000111", -- 10246 FREE #<CONS 0 10247>
 "00000000000000000010100000001000", -- 10247 FREE #<CONS 0 10248>
 "00000000000000000010100000001001", -- 10248 FREE #<CONS 0 10249>
 "00000000000000000010100000001010", -- 10249 FREE #<CONS 0 10250>
 "00000000000000000010100000001011", -- 10250 FREE #<CONS 0 10251>
 "00000000000000000010100000001100", -- 10251 FREE #<CONS 0 10252>
 "00000000000000000010100000001101", -- 10252 FREE #<CONS 0 10253>
 "00000000000000000010100000001110", -- 10253 FREE #<CONS 0 10254>
 "00000000000000000010100000001111", -- 10254 FREE #<CONS 0 10255>
 "00000000000000000010100000010000", -- 10255 FREE #<CONS 0 10256>
 "00000000000000000010100000010001", -- 10256 FREE #<CONS 0 10257>
 "00000000000000000010100000010010", -- 10257 FREE #<CONS 0 10258>
 "00000000000000000010100000010011", -- 10258 FREE #<CONS 0 10259>
 "00000000000000000010100000010100", -- 10259 FREE #<CONS 0 10260>
 "00000000000000000010100000010101", -- 10260 FREE #<CONS 0 10261>
 "00000000000000000010100000010110", -- 10261 FREE #<CONS 0 10262>
 "00000000000000000010100000010111", -- 10262 FREE #<CONS 0 10263>
 "00000000000000000010100000011000", -- 10263 FREE #<CONS 0 10264>
 "00000000000000000010100000011001", -- 10264 FREE #<CONS 0 10265>
 "00000000000000000010100000011010", -- 10265 FREE #<CONS 0 10266>
 "00000000000000000010100000011011", -- 10266 FREE #<CONS 0 10267>
 "00000000000000000010100000011100", -- 10267 FREE #<CONS 0 10268>
 "00000000000000000010100000011101", -- 10268 FREE #<CONS 0 10269>
 "00000000000000000010100000011110", -- 10269 FREE #<CONS 0 10270>
 "00000000000000000010100000011111", -- 10270 FREE #<CONS 0 10271>
 "00000000000000000010100000100000", -- 10271 FREE #<CONS 0 10272>
 "00000000000000000010100000100001", -- 10272 FREE #<CONS 0 10273>
 "00000000000000000010100000100010", -- 10273 FREE #<CONS 0 10274>
 "00000000000000000010100000100011", -- 10274 FREE #<CONS 0 10275>
 "00000000000000000010100000100100", -- 10275 FREE #<CONS 0 10276>
 "00000000000000000010100000100101", -- 10276 FREE #<CONS 0 10277>
 "00000000000000000010100000100110", -- 10277 FREE #<CONS 0 10278>
 "00000000000000000010100000100111", -- 10278 FREE #<CONS 0 10279>
 "00000000000000000010100000101000", -- 10279 FREE #<CONS 0 10280>
 "00000000000000000010100000101001", -- 10280 FREE #<CONS 0 10281>
 "00000000000000000010100000101010", -- 10281 FREE #<CONS 0 10282>
 "00000000000000000010100000101011", -- 10282 FREE #<CONS 0 10283>
 "00000000000000000010100000101100", -- 10283 FREE #<CONS 0 10284>
 "00000000000000000010100000101101", -- 10284 FREE #<CONS 0 10285>
 "00000000000000000010100000101110", -- 10285 FREE #<CONS 0 10286>
 "00000000000000000010100000101111", -- 10286 FREE #<CONS 0 10287>
 "00000000000000000010100000110000", -- 10287 FREE #<CONS 0 10288>
 "00000000000000000010100000110001", -- 10288 FREE #<CONS 0 10289>
 "00000000000000000010100000110010", -- 10289 FREE #<CONS 0 10290>
 "00000000000000000010100000110011", -- 10290 FREE #<CONS 0 10291>
 "00000000000000000010100000110100", -- 10291 FREE #<CONS 0 10292>
 "00000000000000000010100000110101", -- 10292 FREE #<CONS 0 10293>
 "00000000000000000010100000110110", -- 10293 FREE #<CONS 0 10294>
 "00000000000000000010100000110111", -- 10294 FREE #<CONS 0 10295>
 "00000000000000000010100000111000", -- 10295 FREE #<CONS 0 10296>
 "00000000000000000010100000111001", -- 10296 FREE #<CONS 0 10297>
 "00000000000000000010100000111010", -- 10297 FREE #<CONS 0 10298>
 "00000000000000000010100000111011", -- 10298 FREE #<CONS 0 10299>
 "00000000000000000010100000111100", -- 10299 FREE #<CONS 0 10300>
 "00000000000000000010100000111101", -- 10300 FREE #<CONS 0 10301>
 "00000000000000000010100000111110", -- 10301 FREE #<CONS 0 10302>
 "00000000000000000010100000111111", -- 10302 FREE #<CONS 0 10303>
 "00000000000000000010100001000000", -- 10303 FREE #<CONS 0 10304>
 "00000000000000000010100001000001", -- 10304 FREE #<CONS 0 10305>
 "00000000000000000010100001000010", -- 10305 FREE #<CONS 0 10306>
 "00000000000000000010100001000011", -- 10306 FREE #<CONS 0 10307>
 "00000000000000000010100001000100", -- 10307 FREE #<CONS 0 10308>
 "00000000000000000010100001000101", -- 10308 FREE #<CONS 0 10309>
 "00000000000000000010100001000110", -- 10309 FREE #<CONS 0 10310>
 "00000000000000000010100001000111", -- 10310 FREE #<CONS 0 10311>
 "00000000000000000010100001001000", -- 10311 FREE #<CONS 0 10312>
 "00000000000000000010100001001001", -- 10312 FREE #<CONS 0 10313>
 "00000000000000000010100001001010", -- 10313 FREE #<CONS 0 10314>
 "00000000000000000010100001001011", -- 10314 FREE #<CONS 0 10315>
 "00000000000000000010100001001100", -- 10315 FREE #<CONS 0 10316>
 "00000000000000000010100001001101", -- 10316 FREE #<CONS 0 10317>
 "00000000000000000010100001001110", -- 10317 FREE #<CONS 0 10318>
 "00000000000000000010100001001111", -- 10318 FREE #<CONS 0 10319>
 "00000000000000000010100001010000", -- 10319 FREE #<CONS 0 10320>
 "00000000000000000010100001010001", -- 10320 FREE #<CONS 0 10321>
 "00000000000000000010100001010010", -- 10321 FREE #<CONS 0 10322>
 "00000000000000000010100001010011", -- 10322 FREE #<CONS 0 10323>
 "00000000000000000010100001010100", -- 10323 FREE #<CONS 0 10324>
 "00000000000000000010100001010101", -- 10324 FREE #<CONS 0 10325>
 "00000000000000000010100001010110", -- 10325 FREE #<CONS 0 10326>
 "00000000000000000010100001010111", -- 10326 FREE #<CONS 0 10327>
 "00000000000000000010100001011000", -- 10327 FREE #<CONS 0 10328>
 "00000000000000000010100001011001", -- 10328 FREE #<CONS 0 10329>
 "00000000000000000010100001011010", -- 10329 FREE #<CONS 0 10330>
 "00000000000000000010100001011011", -- 10330 FREE #<CONS 0 10331>
 "00000000000000000010100001011100", -- 10331 FREE #<CONS 0 10332>
 "00000000000000000010100001011101", -- 10332 FREE #<CONS 0 10333>
 "00000000000000000010100001011110", -- 10333 FREE #<CONS 0 10334>
 "00000000000000000010100001011111", -- 10334 FREE #<CONS 0 10335>
 "00000000000000000010100001100000", -- 10335 FREE #<CONS 0 10336>
 "00000000000000000010100001100001", -- 10336 FREE #<CONS 0 10337>
 "00000000000000000010100001100010", -- 10337 FREE #<CONS 0 10338>
 "00000000000000000010100001100011", -- 10338 FREE #<CONS 0 10339>
 "00000000000000000010100001100100", -- 10339 FREE #<CONS 0 10340>
 "00000000000000000010100001100101", -- 10340 FREE #<CONS 0 10341>
 "00000000000000000010100001100110", -- 10341 FREE #<CONS 0 10342>
 "00000000000000000010100001100111", -- 10342 FREE #<CONS 0 10343>
 "00000000000000000010100001101000", -- 10343 FREE #<CONS 0 10344>
 "00000000000000000010100001101001", -- 10344 FREE #<CONS 0 10345>
 "00000000000000000010100001101010", -- 10345 FREE #<CONS 0 10346>
 "00000000000000000010100001101011", -- 10346 FREE #<CONS 0 10347>
 "00000000000000000010100001101100", -- 10347 FREE #<CONS 0 10348>
 "00000000000000000010100001101101", -- 10348 FREE #<CONS 0 10349>
 "00000000000000000010100001101110", -- 10349 FREE #<CONS 0 10350>
 "00000000000000000010100001101111", -- 10350 FREE #<CONS 0 10351>
 "00000000000000000010100001110000", -- 10351 FREE #<CONS 0 10352>
 "00000000000000000010100001110001", -- 10352 FREE #<CONS 0 10353>
 "00000000000000000010100001110010", -- 10353 FREE #<CONS 0 10354>
 "00000000000000000010100001110011", -- 10354 FREE #<CONS 0 10355>
 "00000000000000000010100001110100", -- 10355 FREE #<CONS 0 10356>
 "00000000000000000010100001110101", -- 10356 FREE #<CONS 0 10357>
 "00000000000000000010100001110110", -- 10357 FREE #<CONS 0 10358>
 "00000000000000000010100001110111", -- 10358 FREE #<CONS 0 10359>
 "00000000000000000010100001111000", -- 10359 FREE #<CONS 0 10360>
 "00000000000000000010100001111001", -- 10360 FREE #<CONS 0 10361>
 "00000000000000000010100001111010", -- 10361 FREE #<CONS 0 10362>
 "00000000000000000010100001111011", -- 10362 FREE #<CONS 0 10363>
 "00000000000000000010100001111100", -- 10363 FREE #<CONS 0 10364>
 "00000000000000000010100001111101", -- 10364 FREE #<CONS 0 10365>
 "00000000000000000010100001111110", -- 10365 FREE #<CONS 0 10366>
 "00000000000000000010100001111111", -- 10366 FREE #<CONS 0 10367>
 "00000000000000000010100010000000", -- 10367 FREE #<CONS 0 10368>
 "00000000000000000010100010000001", -- 10368 FREE #<CONS 0 10369>
 "00000000000000000010100010000010", -- 10369 FREE #<CONS 0 10370>
 "00000000000000000010100010000011", -- 10370 FREE #<CONS 0 10371>
 "00000000000000000010100010000100", -- 10371 FREE #<CONS 0 10372>
 "00000000000000000010100010000101", -- 10372 FREE #<CONS 0 10373>
 "00000000000000000010100010000110", -- 10373 FREE #<CONS 0 10374>
 "00000000000000000010100010000111", -- 10374 FREE #<CONS 0 10375>
 "00000000000000000010100010001000", -- 10375 FREE #<CONS 0 10376>
 "00000000000000000010100010001001", -- 10376 FREE #<CONS 0 10377>
 "00000000000000000010100010001010", -- 10377 FREE #<CONS 0 10378>
 "00000000000000000010100010001011", -- 10378 FREE #<CONS 0 10379>
 "00000000000000000010100010001100", -- 10379 FREE #<CONS 0 10380>
 "00000000000000000010100010001101", -- 10380 FREE #<CONS 0 10381>
 "00000000000000000010100010001110", -- 10381 FREE #<CONS 0 10382>
 "00000000000000000010100010001111", -- 10382 FREE #<CONS 0 10383>
 "00000000000000000010100010010000", -- 10383 FREE #<CONS 0 10384>
 "00000000000000000010100010010001", -- 10384 FREE #<CONS 0 10385>
 "00000000000000000010100010010010", -- 10385 FREE #<CONS 0 10386>
 "00000000000000000010100010010011", -- 10386 FREE #<CONS 0 10387>
 "00000000000000000010100010010100", -- 10387 FREE #<CONS 0 10388>
 "00000000000000000010100010010101", -- 10388 FREE #<CONS 0 10389>
 "00000000000000000010100010010110", -- 10389 FREE #<CONS 0 10390>
 "00000000000000000010100010010111", -- 10390 FREE #<CONS 0 10391>
 "00000000000000000010100010011000", -- 10391 FREE #<CONS 0 10392>
 "00000000000000000010100010011001", -- 10392 FREE #<CONS 0 10393>
 "00000000000000000010100010011010", -- 10393 FREE #<CONS 0 10394>
 "00000000000000000010100010011011", -- 10394 FREE #<CONS 0 10395>
 "00000000000000000010100010011100", -- 10395 FREE #<CONS 0 10396>
 "00000000000000000010100010011101", -- 10396 FREE #<CONS 0 10397>
 "00000000000000000010100010011110", -- 10397 FREE #<CONS 0 10398>
 "00000000000000000010100010011111", -- 10398 FREE #<CONS 0 10399>
 "00000000000000000010100010100000", -- 10399 FREE #<CONS 0 10400>
 "00000000000000000010100010100001", -- 10400 FREE #<CONS 0 10401>
 "00000000000000000010100010100010", -- 10401 FREE #<CONS 0 10402>
 "00000000000000000010100010100011", -- 10402 FREE #<CONS 0 10403>
 "00000000000000000010100010100100", -- 10403 FREE #<CONS 0 10404>
 "00000000000000000010100010100101", -- 10404 FREE #<CONS 0 10405>
 "00000000000000000010100010100110", -- 10405 FREE #<CONS 0 10406>
 "00000000000000000010100010100111", -- 10406 FREE #<CONS 0 10407>
 "00000000000000000010100010101000", -- 10407 FREE #<CONS 0 10408>
 "00000000000000000010100010101001", -- 10408 FREE #<CONS 0 10409>
 "00000000000000000010100010101010", -- 10409 FREE #<CONS 0 10410>
 "00000000000000000010100010101011", -- 10410 FREE #<CONS 0 10411>
 "00000000000000000010100010101100", -- 10411 FREE #<CONS 0 10412>
 "00000000000000000010100010101101", -- 10412 FREE #<CONS 0 10413>
 "00000000000000000010100010101110", -- 10413 FREE #<CONS 0 10414>
 "00000000000000000010100010101111", -- 10414 FREE #<CONS 0 10415>
 "00000000000000000010100010110000", -- 10415 FREE #<CONS 0 10416>
 "00000000000000000010100010110001", -- 10416 FREE #<CONS 0 10417>
 "00000000000000000010100010110010", -- 10417 FREE #<CONS 0 10418>
 "00000000000000000010100010110011", -- 10418 FREE #<CONS 0 10419>
 "00000000000000000010100010110100", -- 10419 FREE #<CONS 0 10420>
 "00000000000000000010100010110101", -- 10420 FREE #<CONS 0 10421>
 "00000000000000000010100010110110", -- 10421 FREE #<CONS 0 10422>
 "00000000000000000010100010110111", -- 10422 FREE #<CONS 0 10423>
 "00000000000000000010100010111000", -- 10423 FREE #<CONS 0 10424>
 "00000000000000000010100010111001", -- 10424 FREE #<CONS 0 10425>
 "00000000000000000010100010111010", -- 10425 FREE #<CONS 0 10426>
 "00000000000000000010100010111011", -- 10426 FREE #<CONS 0 10427>
 "00000000000000000010100010111100", -- 10427 FREE #<CONS 0 10428>
 "00000000000000000010100010111101", -- 10428 FREE #<CONS 0 10429>
 "00000000000000000010100010111110", -- 10429 FREE #<CONS 0 10430>
 "00000000000000000010100010111111", -- 10430 FREE #<CONS 0 10431>
 "00000000000000000010100011000000", -- 10431 FREE #<CONS 0 10432>
 "00000000000000000010100011000001", -- 10432 FREE #<CONS 0 10433>
 "00000000000000000010100011000010", -- 10433 FREE #<CONS 0 10434>
 "00000000000000000010100011000011", -- 10434 FREE #<CONS 0 10435>
 "00000000000000000010100011000100", -- 10435 FREE #<CONS 0 10436>
 "00000000000000000010100011000101", -- 10436 FREE #<CONS 0 10437>
 "00000000000000000010100011000110", -- 10437 FREE #<CONS 0 10438>
 "00000000000000000010100011000111", -- 10438 FREE #<CONS 0 10439>
 "00000000000000000010100011001000", -- 10439 FREE #<CONS 0 10440>
 "00000000000000000010100011001001", -- 10440 FREE #<CONS 0 10441>
 "00000000000000000010100011001010", -- 10441 FREE #<CONS 0 10442>
 "00000000000000000010100011001011", -- 10442 FREE #<CONS 0 10443>
 "00000000000000000010100011001100", -- 10443 FREE #<CONS 0 10444>
 "00000000000000000010100011001101", -- 10444 FREE #<CONS 0 10445>
 "00000000000000000010100011001110", -- 10445 FREE #<CONS 0 10446>
 "00000000000000000010100011001111", -- 10446 FREE #<CONS 0 10447>
 "00000000000000000010100011010000", -- 10447 FREE #<CONS 0 10448>
 "00000000000000000010100011010001", -- 10448 FREE #<CONS 0 10449>
 "00000000000000000010100011010010", -- 10449 FREE #<CONS 0 10450>
 "00000000000000000010100011010011", -- 10450 FREE #<CONS 0 10451>
 "00000000000000000010100011010100", -- 10451 FREE #<CONS 0 10452>
 "00000000000000000010100011010101", -- 10452 FREE #<CONS 0 10453>
 "00000000000000000010100011010110", -- 10453 FREE #<CONS 0 10454>
 "00000000000000000010100011010111", -- 10454 FREE #<CONS 0 10455>
 "00000000000000000010100011011000", -- 10455 FREE #<CONS 0 10456>
 "00000000000000000010100011011001", -- 10456 FREE #<CONS 0 10457>
 "00000000000000000010100011011010", -- 10457 FREE #<CONS 0 10458>
 "00000000000000000010100011011011", -- 10458 FREE #<CONS 0 10459>
 "00000000000000000010100011011100", -- 10459 FREE #<CONS 0 10460>
 "00000000000000000010100011011101", -- 10460 FREE #<CONS 0 10461>
 "00000000000000000010100011011110", -- 10461 FREE #<CONS 0 10462>
 "00000000000000000010100011011111", -- 10462 FREE #<CONS 0 10463>
 "00000000000000000010100011100000", -- 10463 FREE #<CONS 0 10464>
 "00000000000000000010100011100001", -- 10464 FREE #<CONS 0 10465>
 "00000000000000000010100011100010", -- 10465 FREE #<CONS 0 10466>
 "00000000000000000010100011100011", -- 10466 FREE #<CONS 0 10467>
 "00000000000000000010100011100100", -- 10467 FREE #<CONS 0 10468>
 "00000000000000000010100011100101", -- 10468 FREE #<CONS 0 10469>
 "00000000000000000010100011100110", -- 10469 FREE #<CONS 0 10470>
 "00000000000000000010100011100111", -- 10470 FREE #<CONS 0 10471>
 "00000000000000000010100011101000", -- 10471 FREE #<CONS 0 10472>
 "00000000000000000010100011101001", -- 10472 FREE #<CONS 0 10473>
 "00000000000000000010100011101010", -- 10473 FREE #<CONS 0 10474>
 "00000000000000000010100011101011", -- 10474 FREE #<CONS 0 10475>
 "00000000000000000010100011101100", -- 10475 FREE #<CONS 0 10476>
 "00000000000000000010100011101101", -- 10476 FREE #<CONS 0 10477>
 "00000000000000000010100011101110", -- 10477 FREE #<CONS 0 10478>
 "00000000000000000010100011101111", -- 10478 FREE #<CONS 0 10479>
 "00000000000000000010100011110000", -- 10479 FREE #<CONS 0 10480>
 "00000000000000000010100011110001", -- 10480 FREE #<CONS 0 10481>
 "00000000000000000010100011110010", -- 10481 FREE #<CONS 0 10482>
 "00000000000000000010100011110011", -- 10482 FREE #<CONS 0 10483>
 "00000000000000000010100011110100", -- 10483 FREE #<CONS 0 10484>
 "00000000000000000010100011110101", -- 10484 FREE #<CONS 0 10485>
 "00000000000000000010100011110110", -- 10485 FREE #<CONS 0 10486>
 "00000000000000000010100011110111", -- 10486 FREE #<CONS 0 10487>
 "00000000000000000010100011111000", -- 10487 FREE #<CONS 0 10488>
 "00000000000000000010100011111001", -- 10488 FREE #<CONS 0 10489>
 "00000000000000000010100011111010", -- 10489 FREE #<CONS 0 10490>
 "00000000000000000010100011111011", -- 10490 FREE #<CONS 0 10491>
 "00000000000000000010100011111100", -- 10491 FREE #<CONS 0 10492>
 "00000000000000000010100011111101", -- 10492 FREE #<CONS 0 10493>
 "00000000000000000010100011111110", -- 10493 FREE #<CONS 0 10494>
 "00000000000000000010100011111111", -- 10494 FREE #<CONS 0 10495>
 "00000000000000000010100100000000", -- 10495 FREE #<CONS 0 10496>
 "00000000000000000010100100000001", -- 10496 FREE #<CONS 0 10497>
 "00000000000000000010100100000010", -- 10497 FREE #<CONS 0 10498>
 "00000000000000000010100100000011", -- 10498 FREE #<CONS 0 10499>
 "00000000000000000010100100000100", -- 10499 FREE #<CONS 0 10500>
 "00000000000000000010100100000101", -- 10500 FREE #<CONS 0 10501>
 "00000000000000000010100100000110", -- 10501 FREE #<CONS 0 10502>
 "00000000000000000010100100000111", -- 10502 FREE #<CONS 0 10503>
 "00000000000000000010100100001000", -- 10503 FREE #<CONS 0 10504>
 "00000000000000000010100100001001", -- 10504 FREE #<CONS 0 10505>
 "00000000000000000010100100001010", -- 10505 FREE #<CONS 0 10506>
 "00000000000000000010100100001011", -- 10506 FREE #<CONS 0 10507>
 "00000000000000000010100100001100", -- 10507 FREE #<CONS 0 10508>
 "00000000000000000010100100001101", -- 10508 FREE #<CONS 0 10509>
 "00000000000000000010100100001110", -- 10509 FREE #<CONS 0 10510>
 "00000000000000000010100100001111", -- 10510 FREE #<CONS 0 10511>
 "00000000000000000010100100010000", -- 10511 FREE #<CONS 0 10512>
 "00000000000000000010100100010001", -- 10512 FREE #<CONS 0 10513>
 "00000000000000000010100100010010", -- 10513 FREE #<CONS 0 10514>
 "00000000000000000010100100010011", -- 10514 FREE #<CONS 0 10515>
 "00000000000000000010100100010100", -- 10515 FREE #<CONS 0 10516>
 "00000000000000000010100100010101", -- 10516 FREE #<CONS 0 10517>
 "00000000000000000010100100010110", -- 10517 FREE #<CONS 0 10518>
 "00000000000000000010100100010111", -- 10518 FREE #<CONS 0 10519>
 "00000000000000000010100100011000", -- 10519 FREE #<CONS 0 10520>
 "00000000000000000010100100011001", -- 10520 FREE #<CONS 0 10521>
 "00000000000000000010100100011010", -- 10521 FREE #<CONS 0 10522>
 "00000000000000000010100100011011", -- 10522 FREE #<CONS 0 10523>
 "00000000000000000010100100011100", -- 10523 FREE #<CONS 0 10524>
 "00000000000000000010100100011101", -- 10524 FREE #<CONS 0 10525>
 "00000000000000000010100100011110", -- 10525 FREE #<CONS 0 10526>
 "00000000000000000010100100011111", -- 10526 FREE #<CONS 0 10527>
 "00000000000000000010100100100000", -- 10527 FREE #<CONS 0 10528>
 "00000000000000000010100100100001", -- 10528 FREE #<CONS 0 10529>
 "00000000000000000010100100100010", -- 10529 FREE #<CONS 0 10530>
 "00000000000000000010100100100011", -- 10530 FREE #<CONS 0 10531>
 "00000000000000000010100100100100", -- 10531 FREE #<CONS 0 10532>
 "00000000000000000010100100100101", -- 10532 FREE #<CONS 0 10533>
 "00000000000000000010100100100110", -- 10533 FREE #<CONS 0 10534>
 "00000000000000000010100100100111", -- 10534 FREE #<CONS 0 10535>
 "00000000000000000010100100101000", -- 10535 FREE #<CONS 0 10536>
 "00000000000000000010100100101001", -- 10536 FREE #<CONS 0 10537>
 "00000000000000000010100100101010", -- 10537 FREE #<CONS 0 10538>
 "00000000000000000010100100101011", -- 10538 FREE #<CONS 0 10539>
 "00000000000000000010100100101100", -- 10539 FREE #<CONS 0 10540>
 "00000000000000000010100100101101", -- 10540 FREE #<CONS 0 10541>
 "00000000000000000010100100101110", -- 10541 FREE #<CONS 0 10542>
 "00000000000000000010100100101111", -- 10542 FREE #<CONS 0 10543>
 "00000000000000000010100100110000", -- 10543 FREE #<CONS 0 10544>
 "00000000000000000010100100110001", -- 10544 FREE #<CONS 0 10545>
 "00000000000000000010100100110010", -- 10545 FREE #<CONS 0 10546>
 "00000000000000000010100100110011", -- 10546 FREE #<CONS 0 10547>
 "00000000000000000010100100110100", -- 10547 FREE #<CONS 0 10548>
 "00000000000000000010100100110101", -- 10548 FREE #<CONS 0 10549>
 "00000000000000000010100100110110", -- 10549 FREE #<CONS 0 10550>
 "00000000000000000010100100110111", -- 10550 FREE #<CONS 0 10551>
 "00000000000000000010100100111000", -- 10551 FREE #<CONS 0 10552>
 "00000000000000000010100100111001", -- 10552 FREE #<CONS 0 10553>
 "00000000000000000010100100111010", -- 10553 FREE #<CONS 0 10554>
 "00000000000000000010100100111011", -- 10554 FREE #<CONS 0 10555>
 "00000000000000000010100100111100", -- 10555 FREE #<CONS 0 10556>
 "00000000000000000010100100111101", -- 10556 FREE #<CONS 0 10557>
 "00000000000000000010100100111110", -- 10557 FREE #<CONS 0 10558>
 "00000000000000000010100100111111", -- 10558 FREE #<CONS 0 10559>
 "00000000000000000010100101000000", -- 10559 FREE #<CONS 0 10560>
 "00000000000000000010100101000001", -- 10560 FREE #<CONS 0 10561>
 "00000000000000000010100101000010", -- 10561 FREE #<CONS 0 10562>
 "00000000000000000010100101000011", -- 10562 FREE #<CONS 0 10563>
 "00000000000000000010100101000100", -- 10563 FREE #<CONS 0 10564>
 "00000000000000000010100101000101", -- 10564 FREE #<CONS 0 10565>
 "00000000000000000010100101000110", -- 10565 FREE #<CONS 0 10566>
 "00000000000000000010100101000111", -- 10566 FREE #<CONS 0 10567>
 "00000000000000000010100101001000", -- 10567 FREE #<CONS 0 10568>
 "00000000000000000010100101001001", -- 10568 FREE #<CONS 0 10569>
 "00000000000000000010100101001010", -- 10569 FREE #<CONS 0 10570>
 "00000000000000000010100101001011", -- 10570 FREE #<CONS 0 10571>
 "00000000000000000010100101001100", -- 10571 FREE #<CONS 0 10572>
 "00000000000000000010100101001101", -- 10572 FREE #<CONS 0 10573>
 "00000000000000000010100101001110", -- 10573 FREE #<CONS 0 10574>
 "00000000000000000010100101001111", -- 10574 FREE #<CONS 0 10575>
 "00000000000000000010100101010000", -- 10575 FREE #<CONS 0 10576>
 "00000000000000000010100101010001", -- 10576 FREE #<CONS 0 10577>
 "00000000000000000010100101010010", -- 10577 FREE #<CONS 0 10578>
 "00000000000000000010100101010011", -- 10578 FREE #<CONS 0 10579>
 "00000000000000000010100101010100", -- 10579 FREE #<CONS 0 10580>
 "00000000000000000010100101010101", -- 10580 FREE #<CONS 0 10581>
 "00000000000000000010100101010110", -- 10581 FREE #<CONS 0 10582>
 "00000000000000000010100101010111", -- 10582 FREE #<CONS 0 10583>
 "00000000000000000010100101011000", -- 10583 FREE #<CONS 0 10584>
 "00000000000000000010100101011001", -- 10584 FREE #<CONS 0 10585>
 "00000000000000000010100101011010", -- 10585 FREE #<CONS 0 10586>
 "00000000000000000010100101011011", -- 10586 FREE #<CONS 0 10587>
 "00000000000000000010100101011100", -- 10587 FREE #<CONS 0 10588>
 "00000000000000000010100101011101", -- 10588 FREE #<CONS 0 10589>
 "00000000000000000010100101011110", -- 10589 FREE #<CONS 0 10590>
 "00000000000000000010100101011111", -- 10590 FREE #<CONS 0 10591>
 "00000000000000000010100101100000", -- 10591 FREE #<CONS 0 10592>
 "00000000000000000010100101100001", -- 10592 FREE #<CONS 0 10593>
 "00000000000000000010100101100010", -- 10593 FREE #<CONS 0 10594>
 "00000000000000000010100101100011", -- 10594 FREE #<CONS 0 10595>
 "00000000000000000010100101100100", -- 10595 FREE #<CONS 0 10596>
 "00000000000000000010100101100101", -- 10596 FREE #<CONS 0 10597>
 "00000000000000000010100101100110", -- 10597 FREE #<CONS 0 10598>
 "00000000000000000010100101100111", -- 10598 FREE #<CONS 0 10599>
 "00000000000000000010100101101000", -- 10599 FREE #<CONS 0 10600>
 "00000000000000000010100101101001", -- 10600 FREE #<CONS 0 10601>
 "00000000000000000010100101101010", -- 10601 FREE #<CONS 0 10602>
 "00000000000000000010100101101011", -- 10602 FREE #<CONS 0 10603>
 "00000000000000000010100101101100", -- 10603 FREE #<CONS 0 10604>
 "00000000000000000010100101101101", -- 10604 FREE #<CONS 0 10605>
 "00000000000000000010100101101110", -- 10605 FREE #<CONS 0 10606>
 "00000000000000000010100101101111", -- 10606 FREE #<CONS 0 10607>
 "00000000000000000010100101110000", -- 10607 FREE #<CONS 0 10608>
 "00000000000000000010100101110001", -- 10608 FREE #<CONS 0 10609>
 "00000000000000000010100101110010", -- 10609 FREE #<CONS 0 10610>
 "00000000000000000010100101110011", -- 10610 FREE #<CONS 0 10611>
 "00000000000000000010100101110100", -- 10611 FREE #<CONS 0 10612>
 "00000000000000000010100101110101", -- 10612 FREE #<CONS 0 10613>
 "00000000000000000010100101110110", -- 10613 FREE #<CONS 0 10614>
 "00000000000000000010100101110111", -- 10614 FREE #<CONS 0 10615>
 "00000000000000000010100101111000", -- 10615 FREE #<CONS 0 10616>
 "00000000000000000010100101111001", -- 10616 FREE #<CONS 0 10617>
 "00000000000000000010100101111010", -- 10617 FREE #<CONS 0 10618>
 "00000000000000000010100101111011", -- 10618 FREE #<CONS 0 10619>
 "00000000000000000010100101111100", -- 10619 FREE #<CONS 0 10620>
 "00000000000000000010100101111101", -- 10620 FREE #<CONS 0 10621>
 "00000000000000000010100101111110", -- 10621 FREE #<CONS 0 10622>
 "00000000000000000010100101111111", -- 10622 FREE #<CONS 0 10623>
 "00000000000000000010100110000000", -- 10623 FREE #<CONS 0 10624>
 "00000000000000000010100110000001", -- 10624 FREE #<CONS 0 10625>
 "00000000000000000010100110000010", -- 10625 FREE #<CONS 0 10626>
 "00000000000000000010100110000011", -- 10626 FREE #<CONS 0 10627>
 "00000000000000000010100110000100", -- 10627 FREE #<CONS 0 10628>
 "00000000000000000010100110000101", -- 10628 FREE #<CONS 0 10629>
 "00000000000000000010100110000110", -- 10629 FREE #<CONS 0 10630>
 "00000000000000000010100110000111", -- 10630 FREE #<CONS 0 10631>
 "00000000000000000010100110001000", -- 10631 FREE #<CONS 0 10632>
 "00000000000000000010100110001001", -- 10632 FREE #<CONS 0 10633>
 "00000000000000000010100110001010", -- 10633 FREE #<CONS 0 10634>
 "00000000000000000010100110001011", -- 10634 FREE #<CONS 0 10635>
 "00000000000000000010100110001100", -- 10635 FREE #<CONS 0 10636>
 "00000000000000000010100110001101", -- 10636 FREE #<CONS 0 10637>
 "00000000000000000010100110001110", -- 10637 FREE #<CONS 0 10638>
 "00000000000000000010100110001111", -- 10638 FREE #<CONS 0 10639>
 "00000000000000000010100110010000", -- 10639 FREE #<CONS 0 10640>
 "00000000000000000010100110010001", -- 10640 FREE #<CONS 0 10641>
 "00000000000000000010100110010010", -- 10641 FREE #<CONS 0 10642>
 "00000000000000000010100110010011", -- 10642 FREE #<CONS 0 10643>
 "00000000000000000010100110010100", -- 10643 FREE #<CONS 0 10644>
 "00000000000000000010100110010101", -- 10644 FREE #<CONS 0 10645>
 "00000000000000000010100110010110", -- 10645 FREE #<CONS 0 10646>
 "00000000000000000010100110010111", -- 10646 FREE #<CONS 0 10647>
 "00000000000000000010100110011000", -- 10647 FREE #<CONS 0 10648>
 "00000000000000000010100110011001", -- 10648 FREE #<CONS 0 10649>
 "00000000000000000010100110011010", -- 10649 FREE #<CONS 0 10650>
 "00000000000000000010100110011011", -- 10650 FREE #<CONS 0 10651>
 "00000000000000000010100110011100", -- 10651 FREE #<CONS 0 10652>
 "00000000000000000010100110011101", -- 10652 FREE #<CONS 0 10653>
 "00000000000000000010100110011110", -- 10653 FREE #<CONS 0 10654>
 "00000000000000000010100110011111", -- 10654 FREE #<CONS 0 10655>
 "00000000000000000010100110100000", -- 10655 FREE #<CONS 0 10656>
 "00000000000000000010100110100001", -- 10656 FREE #<CONS 0 10657>
 "00000000000000000010100110100010", -- 10657 FREE #<CONS 0 10658>
 "00000000000000000010100110100011", -- 10658 FREE #<CONS 0 10659>
 "00000000000000000010100110100100", -- 10659 FREE #<CONS 0 10660>
 "00000000000000000010100110100101", -- 10660 FREE #<CONS 0 10661>
 "00000000000000000010100110100110", -- 10661 FREE #<CONS 0 10662>
 "00000000000000000010100110100111", -- 10662 FREE #<CONS 0 10663>
 "00000000000000000010100110101000", -- 10663 FREE #<CONS 0 10664>
 "00000000000000000010100110101001", -- 10664 FREE #<CONS 0 10665>
 "00000000000000000010100110101010", -- 10665 FREE #<CONS 0 10666>
 "00000000000000000010100110101011", -- 10666 FREE #<CONS 0 10667>
 "00000000000000000010100110101100", -- 10667 FREE #<CONS 0 10668>
 "00000000000000000010100110101101", -- 10668 FREE #<CONS 0 10669>
 "00000000000000000010100110101110", -- 10669 FREE #<CONS 0 10670>
 "00000000000000000010100110101111", -- 10670 FREE #<CONS 0 10671>
 "00000000000000000010100110110000", -- 10671 FREE #<CONS 0 10672>
 "00000000000000000010100110110001", -- 10672 FREE #<CONS 0 10673>
 "00000000000000000010100110110010", -- 10673 FREE #<CONS 0 10674>
 "00000000000000000010100110110011", -- 10674 FREE #<CONS 0 10675>
 "00000000000000000010100110110100", -- 10675 FREE #<CONS 0 10676>
 "00000000000000000010100110110101", -- 10676 FREE #<CONS 0 10677>
 "00000000000000000010100110110110", -- 10677 FREE #<CONS 0 10678>
 "00000000000000000010100110110111", -- 10678 FREE #<CONS 0 10679>
 "00000000000000000010100110111000", -- 10679 FREE #<CONS 0 10680>
 "00000000000000000010100110111001", -- 10680 FREE #<CONS 0 10681>
 "00000000000000000010100110111010", -- 10681 FREE #<CONS 0 10682>
 "00000000000000000010100110111011", -- 10682 FREE #<CONS 0 10683>
 "00000000000000000010100110111100", -- 10683 FREE #<CONS 0 10684>
 "00000000000000000010100110111101", -- 10684 FREE #<CONS 0 10685>
 "00000000000000000010100110111110", -- 10685 FREE #<CONS 0 10686>
 "00000000000000000010100110111111", -- 10686 FREE #<CONS 0 10687>
 "00000000000000000010100111000000", -- 10687 FREE #<CONS 0 10688>
 "00000000000000000010100111000001", -- 10688 FREE #<CONS 0 10689>
 "00000000000000000010100111000010", -- 10689 FREE #<CONS 0 10690>
 "00000000000000000010100111000011", -- 10690 FREE #<CONS 0 10691>
 "00000000000000000010100111000100", -- 10691 FREE #<CONS 0 10692>
 "00000000000000000010100111000101", -- 10692 FREE #<CONS 0 10693>
 "00000000000000000010100111000110", -- 10693 FREE #<CONS 0 10694>
 "00000000000000000010100111000111", -- 10694 FREE #<CONS 0 10695>
 "00000000000000000010100111001000", -- 10695 FREE #<CONS 0 10696>
 "00000000000000000010100111001001", -- 10696 FREE #<CONS 0 10697>
 "00000000000000000010100111001010", -- 10697 FREE #<CONS 0 10698>
 "00000000000000000010100111001011", -- 10698 FREE #<CONS 0 10699>
 "00000000000000000010100111001100", -- 10699 FREE #<CONS 0 10700>
 "00000000000000000010100111001101", -- 10700 FREE #<CONS 0 10701>
 "00000000000000000010100111001110", -- 10701 FREE #<CONS 0 10702>
 "00000000000000000010100111001111", -- 10702 FREE #<CONS 0 10703>
 "00000000000000000010100111010000", -- 10703 FREE #<CONS 0 10704>
 "00000000000000000010100111010001", -- 10704 FREE #<CONS 0 10705>
 "00000000000000000010100111010010", -- 10705 FREE #<CONS 0 10706>
 "00000000000000000010100111010011", -- 10706 FREE #<CONS 0 10707>
 "00000000000000000010100111010100", -- 10707 FREE #<CONS 0 10708>
 "00000000000000000010100111010101", -- 10708 FREE #<CONS 0 10709>
 "00000000000000000010100111010110", -- 10709 FREE #<CONS 0 10710>
 "00000000000000000010100111010111", -- 10710 FREE #<CONS 0 10711>
 "00000000000000000010100111011000", -- 10711 FREE #<CONS 0 10712>
 "00000000000000000010100111011001", -- 10712 FREE #<CONS 0 10713>
 "00000000000000000010100111011010", -- 10713 FREE #<CONS 0 10714>
 "00000000000000000010100111011011", -- 10714 FREE #<CONS 0 10715>
 "00000000000000000010100111011100", -- 10715 FREE #<CONS 0 10716>
 "00000000000000000010100111011101", -- 10716 FREE #<CONS 0 10717>
 "00000000000000000010100111011110", -- 10717 FREE #<CONS 0 10718>
 "00000000000000000010100111011111", -- 10718 FREE #<CONS 0 10719>
 "00000000000000000010100111100000", -- 10719 FREE #<CONS 0 10720>
 "00000000000000000010100111100001", -- 10720 FREE #<CONS 0 10721>
 "00000000000000000010100111100010", -- 10721 FREE #<CONS 0 10722>
 "00000000000000000010100111100011", -- 10722 FREE #<CONS 0 10723>
 "00000000000000000010100111100100", -- 10723 FREE #<CONS 0 10724>
 "00000000000000000010100111100101", -- 10724 FREE #<CONS 0 10725>
 "00000000000000000010100111100110", -- 10725 FREE #<CONS 0 10726>
 "00000000000000000010100111100111", -- 10726 FREE #<CONS 0 10727>
 "00000000000000000010100111101000", -- 10727 FREE #<CONS 0 10728>
 "00000000000000000010100111101001", -- 10728 FREE #<CONS 0 10729>
 "00000000000000000010100111101010", -- 10729 FREE #<CONS 0 10730>
 "00000000000000000010100111101011", -- 10730 FREE #<CONS 0 10731>
 "00000000000000000010100111101100", -- 10731 FREE #<CONS 0 10732>
 "00000000000000000010100111101101", -- 10732 FREE #<CONS 0 10733>
 "00000000000000000010100111101110", -- 10733 FREE #<CONS 0 10734>
 "00000000000000000010100111101111", -- 10734 FREE #<CONS 0 10735>
 "00000000000000000010100111110000", -- 10735 FREE #<CONS 0 10736>
 "00000000000000000010100111110001", -- 10736 FREE #<CONS 0 10737>
 "00000000000000000010100111110010", -- 10737 FREE #<CONS 0 10738>
 "00000000000000000010100111110011", -- 10738 FREE #<CONS 0 10739>
 "00000000000000000010100111110100", -- 10739 FREE #<CONS 0 10740>
 "00000000000000000010100111110101", -- 10740 FREE #<CONS 0 10741>
 "00000000000000000010100111110110", -- 10741 FREE #<CONS 0 10742>
 "00000000000000000010100111110111", -- 10742 FREE #<CONS 0 10743>
 "00000000000000000010100111111000", -- 10743 FREE #<CONS 0 10744>
 "00000000000000000010100111111001", -- 10744 FREE #<CONS 0 10745>
 "00000000000000000010100111111010", -- 10745 FREE #<CONS 0 10746>
 "00000000000000000010100111111011", -- 10746 FREE #<CONS 0 10747>
 "00000000000000000010100111111100", -- 10747 FREE #<CONS 0 10748>
 "00000000000000000010100111111101", -- 10748 FREE #<CONS 0 10749>
 "00000000000000000010100111111110", -- 10749 FREE #<CONS 0 10750>
 "00000000000000000010100111111111", -- 10750 FREE #<CONS 0 10751>
 "00000000000000000010101000000000", -- 10751 FREE #<CONS 0 10752>
 "00000000000000000010101000000001", -- 10752 FREE #<CONS 0 10753>
 "00000000000000000010101000000010", -- 10753 FREE #<CONS 0 10754>
 "00000000000000000010101000000011", -- 10754 FREE #<CONS 0 10755>
 "00000000000000000010101000000100", -- 10755 FREE #<CONS 0 10756>
 "00000000000000000010101000000101", -- 10756 FREE #<CONS 0 10757>
 "00000000000000000010101000000110", -- 10757 FREE #<CONS 0 10758>
 "00000000000000000010101000000111", -- 10758 FREE #<CONS 0 10759>
 "00000000000000000010101000001000", -- 10759 FREE #<CONS 0 10760>
 "00000000000000000010101000001001", -- 10760 FREE #<CONS 0 10761>
 "00000000000000000010101000001010", -- 10761 FREE #<CONS 0 10762>
 "00000000000000000010101000001011", -- 10762 FREE #<CONS 0 10763>
 "00000000000000000010101000001100", -- 10763 FREE #<CONS 0 10764>
 "00000000000000000010101000001101", -- 10764 FREE #<CONS 0 10765>
 "00000000000000000010101000001110", -- 10765 FREE #<CONS 0 10766>
 "00000000000000000010101000001111", -- 10766 FREE #<CONS 0 10767>
 "00000000000000000010101000010000", -- 10767 FREE #<CONS 0 10768>
 "00000000000000000010101000010001", -- 10768 FREE #<CONS 0 10769>
 "00000000000000000010101000010010", -- 10769 FREE #<CONS 0 10770>
 "00000000000000000010101000010011", -- 10770 FREE #<CONS 0 10771>
 "00000000000000000010101000010100", -- 10771 FREE #<CONS 0 10772>
 "00000000000000000010101000010101", -- 10772 FREE #<CONS 0 10773>
 "00000000000000000010101000010110", -- 10773 FREE #<CONS 0 10774>
 "00000000000000000010101000010111", -- 10774 FREE #<CONS 0 10775>
 "00000000000000000010101000011000", -- 10775 FREE #<CONS 0 10776>
 "00000000000000000010101000011001", -- 10776 FREE #<CONS 0 10777>
 "00000000000000000010101000011010", -- 10777 FREE #<CONS 0 10778>
 "00000000000000000010101000011011", -- 10778 FREE #<CONS 0 10779>
 "00000000000000000010101000011100", -- 10779 FREE #<CONS 0 10780>
 "00000000000000000010101000011101", -- 10780 FREE #<CONS 0 10781>
 "00000000000000000010101000011110", -- 10781 FREE #<CONS 0 10782>
 "00000000000000000010101000011111", -- 10782 FREE #<CONS 0 10783>
 "00000000000000000010101000100000", -- 10783 FREE #<CONS 0 10784>
 "00000000000000000010101000100001", -- 10784 FREE #<CONS 0 10785>
 "00000000000000000010101000100010", -- 10785 FREE #<CONS 0 10786>
 "00000000000000000010101000100011", -- 10786 FREE #<CONS 0 10787>
 "00000000000000000010101000100100", -- 10787 FREE #<CONS 0 10788>
 "00000000000000000010101000100101", -- 10788 FREE #<CONS 0 10789>
 "00000000000000000010101000100110", -- 10789 FREE #<CONS 0 10790>
 "00000000000000000010101000100111", -- 10790 FREE #<CONS 0 10791>
 "00000000000000000010101000101000", -- 10791 FREE #<CONS 0 10792>
 "00000000000000000010101000101001", -- 10792 FREE #<CONS 0 10793>
 "00000000000000000010101000101010", -- 10793 FREE #<CONS 0 10794>
 "00000000000000000010101000101011", -- 10794 FREE #<CONS 0 10795>
 "00000000000000000010101000101100", -- 10795 FREE #<CONS 0 10796>
 "00000000000000000010101000101101", -- 10796 FREE #<CONS 0 10797>
 "00000000000000000010101000101110", -- 10797 FREE #<CONS 0 10798>
 "00000000000000000010101000101111", -- 10798 FREE #<CONS 0 10799>
 "00000000000000000010101000110000", -- 10799 FREE #<CONS 0 10800>
 "00000000000000000010101000110001", -- 10800 FREE #<CONS 0 10801>
 "00000000000000000010101000110010", -- 10801 FREE #<CONS 0 10802>
 "00000000000000000010101000110011", -- 10802 FREE #<CONS 0 10803>
 "00000000000000000010101000110100", -- 10803 FREE #<CONS 0 10804>
 "00000000000000000010101000110101", -- 10804 FREE #<CONS 0 10805>
 "00000000000000000010101000110110", -- 10805 FREE #<CONS 0 10806>
 "00000000000000000010101000110111", -- 10806 FREE #<CONS 0 10807>
 "00000000000000000010101000111000", -- 10807 FREE #<CONS 0 10808>
 "00000000000000000010101000111001", -- 10808 FREE #<CONS 0 10809>
 "00000000000000000010101000111010", -- 10809 FREE #<CONS 0 10810>
 "00000000000000000010101000111011", -- 10810 FREE #<CONS 0 10811>
 "00000000000000000010101000111100", -- 10811 FREE #<CONS 0 10812>
 "00000000000000000010101000111101", -- 10812 FREE #<CONS 0 10813>
 "00000000000000000010101000111110", -- 10813 FREE #<CONS 0 10814>
 "00000000000000000010101000111111", -- 10814 FREE #<CONS 0 10815>
 "00000000000000000010101001000000", -- 10815 FREE #<CONS 0 10816>
 "00000000000000000010101001000001", -- 10816 FREE #<CONS 0 10817>
 "00000000000000000010101001000010", -- 10817 FREE #<CONS 0 10818>
 "00000000000000000010101001000011", -- 10818 FREE #<CONS 0 10819>
 "00000000000000000010101001000100", -- 10819 FREE #<CONS 0 10820>
 "00000000000000000010101001000101", -- 10820 FREE #<CONS 0 10821>
 "00000000000000000010101001000110", -- 10821 FREE #<CONS 0 10822>
 "00000000000000000010101001000111", -- 10822 FREE #<CONS 0 10823>
 "00000000000000000010101001001000", -- 10823 FREE #<CONS 0 10824>
 "00000000000000000010101001001001", -- 10824 FREE #<CONS 0 10825>
 "00000000000000000010101001001010", -- 10825 FREE #<CONS 0 10826>
 "00000000000000000010101001001011", -- 10826 FREE #<CONS 0 10827>
 "00000000000000000010101001001100", -- 10827 FREE #<CONS 0 10828>
 "00000000000000000010101001001101", -- 10828 FREE #<CONS 0 10829>
 "00000000000000000010101001001110", -- 10829 FREE #<CONS 0 10830>
 "00000000000000000010101001001111", -- 10830 FREE #<CONS 0 10831>
 "00000000000000000010101001010000", -- 10831 FREE #<CONS 0 10832>
 "00000000000000000010101001010001", -- 10832 FREE #<CONS 0 10833>
 "00000000000000000010101001010010", -- 10833 FREE #<CONS 0 10834>
 "00000000000000000010101001010011", -- 10834 FREE #<CONS 0 10835>
 "00000000000000000010101001010100", -- 10835 FREE #<CONS 0 10836>
 "00000000000000000010101001010101", -- 10836 FREE #<CONS 0 10837>
 "00000000000000000010101001010110", -- 10837 FREE #<CONS 0 10838>
 "00000000000000000010101001010111", -- 10838 FREE #<CONS 0 10839>
 "00000000000000000010101001011000", -- 10839 FREE #<CONS 0 10840>
 "00000000000000000010101001011001", -- 10840 FREE #<CONS 0 10841>
 "00000000000000000010101001011010", -- 10841 FREE #<CONS 0 10842>
 "00000000000000000010101001011011", -- 10842 FREE #<CONS 0 10843>
 "00000000000000000010101001011100", -- 10843 FREE #<CONS 0 10844>
 "00000000000000000010101001011101", -- 10844 FREE #<CONS 0 10845>
 "00000000000000000010101001011110", -- 10845 FREE #<CONS 0 10846>
 "00000000000000000010101001011111", -- 10846 FREE #<CONS 0 10847>
 "00000000000000000010101001100000", -- 10847 FREE #<CONS 0 10848>
 "00000000000000000010101001100001", -- 10848 FREE #<CONS 0 10849>
 "00000000000000000010101001100010", -- 10849 FREE #<CONS 0 10850>
 "00000000000000000010101001100011", -- 10850 FREE #<CONS 0 10851>
 "00000000000000000010101001100100", -- 10851 FREE #<CONS 0 10852>
 "00000000000000000010101001100101", -- 10852 FREE #<CONS 0 10853>
 "00000000000000000010101001100110", -- 10853 FREE #<CONS 0 10854>
 "00000000000000000010101001100111", -- 10854 FREE #<CONS 0 10855>
 "00000000000000000010101001101000", -- 10855 FREE #<CONS 0 10856>
 "00000000000000000010101001101001", -- 10856 FREE #<CONS 0 10857>
 "00000000000000000010101001101010", -- 10857 FREE #<CONS 0 10858>
 "00000000000000000010101001101011", -- 10858 FREE #<CONS 0 10859>
 "00000000000000000010101001101100", -- 10859 FREE #<CONS 0 10860>
 "00000000000000000010101001101101", -- 10860 FREE #<CONS 0 10861>
 "00000000000000000010101001101110", -- 10861 FREE #<CONS 0 10862>
 "00000000000000000010101001101111", -- 10862 FREE #<CONS 0 10863>
 "00000000000000000010101001110000", -- 10863 FREE #<CONS 0 10864>
 "00000000000000000010101001110001", -- 10864 FREE #<CONS 0 10865>
 "00000000000000000010101001110010", -- 10865 FREE #<CONS 0 10866>
 "00000000000000000010101001110011", -- 10866 FREE #<CONS 0 10867>
 "00000000000000000010101001110100", -- 10867 FREE #<CONS 0 10868>
 "00000000000000000010101001110101", -- 10868 FREE #<CONS 0 10869>
 "00000000000000000010101001110110", -- 10869 FREE #<CONS 0 10870>
 "00000000000000000010101001110111", -- 10870 FREE #<CONS 0 10871>
 "00000000000000000010101001111000", -- 10871 FREE #<CONS 0 10872>
 "00000000000000000010101001111001", -- 10872 FREE #<CONS 0 10873>
 "00000000000000000010101001111010", -- 10873 FREE #<CONS 0 10874>
 "00000000000000000010101001111011", -- 10874 FREE #<CONS 0 10875>
 "00000000000000000010101001111100", -- 10875 FREE #<CONS 0 10876>
 "00000000000000000010101001111101", -- 10876 FREE #<CONS 0 10877>
 "00000000000000000010101001111110", -- 10877 FREE #<CONS 0 10878>
 "00000000000000000010101001111111", -- 10878 FREE #<CONS 0 10879>
 "00000000000000000010101010000000", -- 10879 FREE #<CONS 0 10880>
 "00000000000000000010101010000001", -- 10880 FREE #<CONS 0 10881>
 "00000000000000000010101010000010", -- 10881 FREE #<CONS 0 10882>
 "00000000000000000010101010000011", -- 10882 FREE #<CONS 0 10883>
 "00000000000000000010101010000100", -- 10883 FREE #<CONS 0 10884>
 "00000000000000000010101010000101", -- 10884 FREE #<CONS 0 10885>
 "00000000000000000010101010000110", -- 10885 FREE #<CONS 0 10886>
 "00000000000000000010101010000111", -- 10886 FREE #<CONS 0 10887>
 "00000000000000000010101010001000", -- 10887 FREE #<CONS 0 10888>
 "00000000000000000010101010001001", -- 10888 FREE #<CONS 0 10889>
 "00000000000000000010101010001010", -- 10889 FREE #<CONS 0 10890>
 "00000000000000000010101010001011", -- 10890 FREE #<CONS 0 10891>
 "00000000000000000010101010001100", -- 10891 FREE #<CONS 0 10892>
 "00000000000000000010101010001101", -- 10892 FREE #<CONS 0 10893>
 "00000000000000000010101010001110", -- 10893 FREE #<CONS 0 10894>
 "00000000000000000010101010001111", -- 10894 FREE #<CONS 0 10895>
 "00000000000000000010101010010000", -- 10895 FREE #<CONS 0 10896>
 "00000000000000000010101010010001", -- 10896 FREE #<CONS 0 10897>
 "00000000000000000010101010010010", -- 10897 FREE #<CONS 0 10898>
 "00000000000000000010101010010011", -- 10898 FREE #<CONS 0 10899>
 "00000000000000000010101010010100", -- 10899 FREE #<CONS 0 10900>
 "00000000000000000010101010010101", -- 10900 FREE #<CONS 0 10901>
 "00000000000000000010101010010110", -- 10901 FREE #<CONS 0 10902>
 "00000000000000000010101010010111", -- 10902 FREE #<CONS 0 10903>
 "00000000000000000010101010011000", -- 10903 FREE #<CONS 0 10904>
 "00000000000000000010101010011001", -- 10904 FREE #<CONS 0 10905>
 "00000000000000000010101010011010", -- 10905 FREE #<CONS 0 10906>
 "00000000000000000010101010011011", -- 10906 FREE #<CONS 0 10907>
 "00000000000000000010101010011100", -- 10907 FREE #<CONS 0 10908>
 "00000000000000000010101010011101", -- 10908 FREE #<CONS 0 10909>
 "00000000000000000010101010011110", -- 10909 FREE #<CONS 0 10910>
 "00000000000000000010101010011111", -- 10910 FREE #<CONS 0 10911>
 "00000000000000000010101010100000", -- 10911 FREE #<CONS 0 10912>
 "00000000000000000010101010100001", -- 10912 FREE #<CONS 0 10913>
 "00000000000000000010101010100010", -- 10913 FREE #<CONS 0 10914>
 "00000000000000000010101010100011", -- 10914 FREE #<CONS 0 10915>
 "00000000000000000010101010100100", -- 10915 FREE #<CONS 0 10916>
 "00000000000000000010101010100101", -- 10916 FREE #<CONS 0 10917>
 "00000000000000000010101010100110", -- 10917 FREE #<CONS 0 10918>
 "00000000000000000010101010100111", -- 10918 FREE #<CONS 0 10919>
 "00000000000000000010101010101000", -- 10919 FREE #<CONS 0 10920>
 "00000000000000000010101010101001", -- 10920 FREE #<CONS 0 10921>
 "00000000000000000010101010101010", -- 10921 FREE #<CONS 0 10922>
 "00000000000000000010101010101011", -- 10922 FREE #<CONS 0 10923>
 "00000000000000000010101010101100", -- 10923 FREE #<CONS 0 10924>
 "00000000000000000010101010101101", -- 10924 FREE #<CONS 0 10925>
 "00000000000000000010101010101110", -- 10925 FREE #<CONS 0 10926>
 "00000000000000000010101010101111", -- 10926 FREE #<CONS 0 10927>
 "00000000000000000010101010110000", -- 10927 FREE #<CONS 0 10928>
 "00000000000000000010101010110001", -- 10928 FREE #<CONS 0 10929>
 "00000000000000000010101010110010", -- 10929 FREE #<CONS 0 10930>
 "00000000000000000010101010110011", -- 10930 FREE #<CONS 0 10931>
 "00000000000000000010101010110100", -- 10931 FREE #<CONS 0 10932>
 "00000000000000000010101010110101", -- 10932 FREE #<CONS 0 10933>
 "00000000000000000010101010110110", -- 10933 FREE #<CONS 0 10934>
 "00000000000000000010101010110111", -- 10934 FREE #<CONS 0 10935>
 "00000000000000000010101010111000", -- 10935 FREE #<CONS 0 10936>
 "00000000000000000010101010111001", -- 10936 FREE #<CONS 0 10937>
 "00000000000000000010101010111010", -- 10937 FREE #<CONS 0 10938>
 "00000000000000000010101010111011", -- 10938 FREE #<CONS 0 10939>
 "00000000000000000010101010111100", -- 10939 FREE #<CONS 0 10940>
 "00000000000000000010101010111101", -- 10940 FREE #<CONS 0 10941>
 "00000000000000000010101010111110", -- 10941 FREE #<CONS 0 10942>
 "00000000000000000010101010111111", -- 10942 FREE #<CONS 0 10943>
 "00000000000000000010101011000000", -- 10943 FREE #<CONS 0 10944>
 "00000000000000000010101011000001", -- 10944 FREE #<CONS 0 10945>
 "00000000000000000010101011000010", -- 10945 FREE #<CONS 0 10946>
 "00000000000000000010101011000011", -- 10946 FREE #<CONS 0 10947>
 "00000000000000000010101011000100", -- 10947 FREE #<CONS 0 10948>
 "00000000000000000010101011000101", -- 10948 FREE #<CONS 0 10949>
 "00000000000000000010101011000110", -- 10949 FREE #<CONS 0 10950>
 "00000000000000000010101011000111", -- 10950 FREE #<CONS 0 10951>
 "00000000000000000010101011001000", -- 10951 FREE #<CONS 0 10952>
 "00000000000000000010101011001001", -- 10952 FREE #<CONS 0 10953>
 "00000000000000000010101011001010", -- 10953 FREE #<CONS 0 10954>
 "00000000000000000010101011001011", -- 10954 FREE #<CONS 0 10955>
 "00000000000000000010101011001100", -- 10955 FREE #<CONS 0 10956>
 "00000000000000000010101011001101", -- 10956 FREE #<CONS 0 10957>
 "00000000000000000010101011001110", -- 10957 FREE #<CONS 0 10958>
 "00000000000000000010101011001111", -- 10958 FREE #<CONS 0 10959>
 "00000000000000000010101011010000", -- 10959 FREE #<CONS 0 10960>
 "00000000000000000010101011010001", -- 10960 FREE #<CONS 0 10961>
 "00000000000000000010101011010010", -- 10961 FREE #<CONS 0 10962>
 "00000000000000000010101011010011", -- 10962 FREE #<CONS 0 10963>
 "00000000000000000010101011010100", -- 10963 FREE #<CONS 0 10964>
 "00000000000000000010101011010101", -- 10964 FREE #<CONS 0 10965>
 "00000000000000000010101011010110", -- 10965 FREE #<CONS 0 10966>
 "00000000000000000010101011010111", -- 10966 FREE #<CONS 0 10967>
 "00000000000000000010101011011000", -- 10967 FREE #<CONS 0 10968>
 "00000000000000000010101011011001", -- 10968 FREE #<CONS 0 10969>
 "00000000000000000010101011011010", -- 10969 FREE #<CONS 0 10970>
 "00000000000000000010101011011011", -- 10970 FREE #<CONS 0 10971>
 "00000000000000000010101011011100", -- 10971 FREE #<CONS 0 10972>
 "00000000000000000010101011011101", -- 10972 FREE #<CONS 0 10973>
 "00000000000000000010101011011110", -- 10973 FREE #<CONS 0 10974>
 "00000000000000000010101011011111", -- 10974 FREE #<CONS 0 10975>
 "00000000000000000010101011100000", -- 10975 FREE #<CONS 0 10976>
 "00000000000000000010101011100001", -- 10976 FREE #<CONS 0 10977>
 "00000000000000000010101011100010", -- 10977 FREE #<CONS 0 10978>
 "00000000000000000010101011100011", -- 10978 FREE #<CONS 0 10979>
 "00000000000000000010101011100100", -- 10979 FREE #<CONS 0 10980>
 "00000000000000000010101011100101", -- 10980 FREE #<CONS 0 10981>
 "00000000000000000010101011100110", -- 10981 FREE #<CONS 0 10982>
 "00000000000000000010101011100111", -- 10982 FREE #<CONS 0 10983>
 "00000000000000000010101011101000", -- 10983 FREE #<CONS 0 10984>
 "00000000000000000010101011101001", -- 10984 FREE #<CONS 0 10985>
 "00000000000000000010101011101010", -- 10985 FREE #<CONS 0 10986>
 "00000000000000000010101011101011", -- 10986 FREE #<CONS 0 10987>
 "00000000000000000010101011101100", -- 10987 FREE #<CONS 0 10988>
 "00000000000000000010101011101101", -- 10988 FREE #<CONS 0 10989>
 "00000000000000000010101011101110", -- 10989 FREE #<CONS 0 10990>
 "00000000000000000010101011101111", -- 10990 FREE #<CONS 0 10991>
 "00000000000000000010101011110000", -- 10991 FREE #<CONS 0 10992>
 "00000000000000000010101011110001", -- 10992 FREE #<CONS 0 10993>
 "00000000000000000010101011110010", -- 10993 FREE #<CONS 0 10994>
 "00000000000000000010101011110011", -- 10994 FREE #<CONS 0 10995>
 "00000000000000000010101011110100", -- 10995 FREE #<CONS 0 10996>
 "00000000000000000010101011110101", -- 10996 FREE #<CONS 0 10997>
 "00000000000000000010101011110110", -- 10997 FREE #<CONS 0 10998>
 "00000000000000000010101011110111", -- 10998 FREE #<CONS 0 10999>
 "00000000000000000010101011111000", -- 10999 FREE #<CONS 0 11000>
 "00000000000000000010101011111001", -- 11000 FREE #<CONS 0 11001>
 "00000000000000000010101011111010", -- 11001 FREE #<CONS 0 11002>
 "00000000000000000010101011111011", -- 11002 FREE #<CONS 0 11003>
 "00000000000000000010101011111100", -- 11003 FREE #<CONS 0 11004>
 "00000000000000000010101011111101", -- 11004 FREE #<CONS 0 11005>
 "00000000000000000010101011111110", -- 11005 FREE #<CONS 0 11006>
 "00000000000000000010101011111111", -- 11006 FREE #<CONS 0 11007>
 "00000000000000000010101100000000", -- 11007 FREE #<CONS 0 11008>
 "00000000000000000010101100000001", -- 11008 FREE #<CONS 0 11009>
 "00000000000000000010101100000010", -- 11009 FREE #<CONS 0 11010>
 "00000000000000000010101100000011", -- 11010 FREE #<CONS 0 11011>
 "00000000000000000010101100000100", -- 11011 FREE #<CONS 0 11012>
 "00000000000000000010101100000101", -- 11012 FREE #<CONS 0 11013>
 "00000000000000000010101100000110", -- 11013 FREE #<CONS 0 11014>
 "00000000000000000010101100000111", -- 11014 FREE #<CONS 0 11015>
 "00000000000000000010101100001000", -- 11015 FREE #<CONS 0 11016>
 "00000000000000000010101100001001", -- 11016 FREE #<CONS 0 11017>
 "00000000000000000010101100001010", -- 11017 FREE #<CONS 0 11018>
 "00000000000000000010101100001011", -- 11018 FREE #<CONS 0 11019>
 "00000000000000000010101100001100", -- 11019 FREE #<CONS 0 11020>
 "00000000000000000010101100001101", -- 11020 FREE #<CONS 0 11021>
 "00000000000000000010101100001110", -- 11021 FREE #<CONS 0 11022>
 "00000000000000000010101100001111", -- 11022 FREE #<CONS 0 11023>
 "00000000000000000010101100010000", -- 11023 FREE #<CONS 0 11024>
 "00000000000000000010101100010001", -- 11024 FREE #<CONS 0 11025>
 "00000000000000000010101100010010", -- 11025 FREE #<CONS 0 11026>
 "00000000000000000010101100010011", -- 11026 FREE #<CONS 0 11027>
 "00000000000000000010101100010100", -- 11027 FREE #<CONS 0 11028>
 "00000000000000000010101100010101", -- 11028 FREE #<CONS 0 11029>
 "00000000000000000010101100010110", -- 11029 FREE #<CONS 0 11030>
 "00000000000000000010101100010111", -- 11030 FREE #<CONS 0 11031>
 "00000000000000000010101100011000", -- 11031 FREE #<CONS 0 11032>
 "00000000000000000010101100011001", -- 11032 FREE #<CONS 0 11033>
 "00000000000000000010101100011010", -- 11033 FREE #<CONS 0 11034>
 "00000000000000000010101100011011", -- 11034 FREE #<CONS 0 11035>
 "00000000000000000010101100011100", -- 11035 FREE #<CONS 0 11036>
 "00000000000000000010101100011101", -- 11036 FREE #<CONS 0 11037>
 "00000000000000000010101100011110", -- 11037 FREE #<CONS 0 11038>
 "00000000000000000010101100011111", -- 11038 FREE #<CONS 0 11039>
 "00000000000000000010101100100000", -- 11039 FREE #<CONS 0 11040>
 "00000000000000000010101100100001", -- 11040 FREE #<CONS 0 11041>
 "00000000000000000010101100100010", -- 11041 FREE #<CONS 0 11042>
 "00000000000000000010101100100011", -- 11042 FREE #<CONS 0 11043>
 "00000000000000000010101100100100", -- 11043 FREE #<CONS 0 11044>
 "00000000000000000010101100100101", -- 11044 FREE #<CONS 0 11045>
 "00000000000000000010101100100110", -- 11045 FREE #<CONS 0 11046>
 "00000000000000000010101100100111", -- 11046 FREE #<CONS 0 11047>
 "00000000000000000010101100101000", -- 11047 FREE #<CONS 0 11048>
 "00000000000000000010101100101001", -- 11048 FREE #<CONS 0 11049>
 "00000000000000000010101100101010", -- 11049 FREE #<CONS 0 11050>
 "00000000000000000010101100101011", -- 11050 FREE #<CONS 0 11051>
 "00000000000000000010101100101100", -- 11051 FREE #<CONS 0 11052>
 "00000000000000000010101100101101", -- 11052 FREE #<CONS 0 11053>
 "00000000000000000010101100101110", -- 11053 FREE #<CONS 0 11054>
 "00000000000000000010101100101111", -- 11054 FREE #<CONS 0 11055>
 "00000000000000000010101100110000", -- 11055 FREE #<CONS 0 11056>
 "00000000000000000010101100110001", -- 11056 FREE #<CONS 0 11057>
 "00000000000000000010101100110010", -- 11057 FREE #<CONS 0 11058>
 "00000000000000000010101100110011", -- 11058 FREE #<CONS 0 11059>
 "00000000000000000010101100110100", -- 11059 FREE #<CONS 0 11060>
 "00000000000000000010101100110101", -- 11060 FREE #<CONS 0 11061>
 "00000000000000000010101100110110", -- 11061 FREE #<CONS 0 11062>
 "00000000000000000010101100110111", -- 11062 FREE #<CONS 0 11063>
 "00000000000000000010101100111000", -- 11063 FREE #<CONS 0 11064>
 "00000000000000000010101100111001", -- 11064 FREE #<CONS 0 11065>
 "00000000000000000010101100111010", -- 11065 FREE #<CONS 0 11066>
 "00000000000000000010101100111011", -- 11066 FREE #<CONS 0 11067>
 "00000000000000000010101100111100", -- 11067 FREE #<CONS 0 11068>
 "00000000000000000010101100111101", -- 11068 FREE #<CONS 0 11069>
 "00000000000000000010101100111110", -- 11069 FREE #<CONS 0 11070>
 "00000000000000000010101100111111", -- 11070 FREE #<CONS 0 11071>
 "00000000000000000010101101000000", -- 11071 FREE #<CONS 0 11072>
 "00000000000000000010101101000001", -- 11072 FREE #<CONS 0 11073>
 "00000000000000000010101101000010", -- 11073 FREE #<CONS 0 11074>
 "00000000000000000010101101000011", -- 11074 FREE #<CONS 0 11075>
 "00000000000000000010101101000100", -- 11075 FREE #<CONS 0 11076>
 "00000000000000000010101101000101", -- 11076 FREE #<CONS 0 11077>
 "00000000000000000010101101000110", -- 11077 FREE #<CONS 0 11078>
 "00000000000000000010101101000111", -- 11078 FREE #<CONS 0 11079>
 "00000000000000000010101101001000", -- 11079 FREE #<CONS 0 11080>
 "00000000000000000010101101001001", -- 11080 FREE #<CONS 0 11081>
 "00000000000000000010101101001010", -- 11081 FREE #<CONS 0 11082>
 "00000000000000000010101101001011", -- 11082 FREE #<CONS 0 11083>
 "00000000000000000010101101001100", -- 11083 FREE #<CONS 0 11084>
 "00000000000000000010101101001101", -- 11084 FREE #<CONS 0 11085>
 "00000000000000000010101101001110", -- 11085 FREE #<CONS 0 11086>
 "00000000000000000010101101001111", -- 11086 FREE #<CONS 0 11087>
 "00000000000000000010101101010000", -- 11087 FREE #<CONS 0 11088>
 "00000000000000000010101101010001", -- 11088 FREE #<CONS 0 11089>
 "00000000000000000010101101010010", -- 11089 FREE #<CONS 0 11090>
 "00000000000000000010101101010011", -- 11090 FREE #<CONS 0 11091>
 "00000000000000000010101101010100", -- 11091 FREE #<CONS 0 11092>
 "00000000000000000010101101010101", -- 11092 FREE #<CONS 0 11093>
 "00000000000000000010101101010110", -- 11093 FREE #<CONS 0 11094>
 "00000000000000000010101101010111", -- 11094 FREE #<CONS 0 11095>
 "00000000000000000010101101011000", -- 11095 FREE #<CONS 0 11096>
 "00000000000000000010101101011001", -- 11096 FREE #<CONS 0 11097>
 "00000000000000000010101101011010", -- 11097 FREE #<CONS 0 11098>
 "00000000000000000010101101011011", -- 11098 FREE #<CONS 0 11099>
 "00000000000000000010101101011100", -- 11099 FREE #<CONS 0 11100>
 "00000000000000000010101101011101", -- 11100 FREE #<CONS 0 11101>
 "00000000000000000010101101011110", -- 11101 FREE #<CONS 0 11102>
 "00000000000000000010101101011111", -- 11102 FREE #<CONS 0 11103>
 "00000000000000000010101101100000", -- 11103 FREE #<CONS 0 11104>
 "00000000000000000010101101100001", -- 11104 FREE #<CONS 0 11105>
 "00000000000000000010101101100010", -- 11105 FREE #<CONS 0 11106>
 "00000000000000000010101101100011", -- 11106 FREE #<CONS 0 11107>
 "00000000000000000010101101100100", -- 11107 FREE #<CONS 0 11108>
 "00000000000000000010101101100101", -- 11108 FREE #<CONS 0 11109>
 "00000000000000000010101101100110", -- 11109 FREE #<CONS 0 11110>
 "00000000000000000010101101100111", -- 11110 FREE #<CONS 0 11111>
 "00000000000000000010101101101000", -- 11111 FREE #<CONS 0 11112>
 "00000000000000000010101101101001", -- 11112 FREE #<CONS 0 11113>
 "00000000000000000010101101101010", -- 11113 FREE #<CONS 0 11114>
 "00000000000000000010101101101011", -- 11114 FREE #<CONS 0 11115>
 "00000000000000000010101101101100", -- 11115 FREE #<CONS 0 11116>
 "00000000000000000010101101101101", -- 11116 FREE #<CONS 0 11117>
 "00000000000000000010101101101110", -- 11117 FREE #<CONS 0 11118>
 "00000000000000000010101101101111", -- 11118 FREE #<CONS 0 11119>
 "00000000000000000010101101110000", -- 11119 FREE #<CONS 0 11120>
 "00000000000000000010101101110001", -- 11120 FREE #<CONS 0 11121>
 "00000000000000000010101101110010", -- 11121 FREE #<CONS 0 11122>
 "00000000000000000010101101110011", -- 11122 FREE #<CONS 0 11123>
 "00000000000000000010101101110100", -- 11123 FREE #<CONS 0 11124>
 "00000000000000000010101101110101", -- 11124 FREE #<CONS 0 11125>
 "00000000000000000010101101110110", -- 11125 FREE #<CONS 0 11126>
 "00000000000000000010101101110111", -- 11126 FREE #<CONS 0 11127>
 "00000000000000000010101101111000", -- 11127 FREE #<CONS 0 11128>
 "00000000000000000010101101111001", -- 11128 FREE #<CONS 0 11129>
 "00000000000000000010101101111010", -- 11129 FREE #<CONS 0 11130>
 "00000000000000000010101101111011", -- 11130 FREE #<CONS 0 11131>
 "00000000000000000010101101111100", -- 11131 FREE #<CONS 0 11132>
 "00000000000000000010101101111101", -- 11132 FREE #<CONS 0 11133>
 "00000000000000000010101101111110", -- 11133 FREE #<CONS 0 11134>
 "00000000000000000010101101111111", -- 11134 FREE #<CONS 0 11135>
 "00000000000000000010101110000000", -- 11135 FREE #<CONS 0 11136>
 "00000000000000000010101110000001", -- 11136 FREE #<CONS 0 11137>
 "00000000000000000010101110000010", -- 11137 FREE #<CONS 0 11138>
 "00000000000000000010101110000011", -- 11138 FREE #<CONS 0 11139>
 "00000000000000000010101110000100", -- 11139 FREE #<CONS 0 11140>
 "00000000000000000010101110000101", -- 11140 FREE #<CONS 0 11141>
 "00000000000000000010101110000110", -- 11141 FREE #<CONS 0 11142>
 "00000000000000000010101110000111", -- 11142 FREE #<CONS 0 11143>
 "00000000000000000010101110001000", -- 11143 FREE #<CONS 0 11144>
 "00000000000000000010101110001001", -- 11144 FREE #<CONS 0 11145>
 "00000000000000000010101110001010", -- 11145 FREE #<CONS 0 11146>
 "00000000000000000010101110001011", -- 11146 FREE #<CONS 0 11147>
 "00000000000000000010101110001100", -- 11147 FREE #<CONS 0 11148>
 "00000000000000000010101110001101", -- 11148 FREE #<CONS 0 11149>
 "00000000000000000010101110001110", -- 11149 FREE #<CONS 0 11150>
 "00000000000000000010101110001111", -- 11150 FREE #<CONS 0 11151>
 "00000000000000000010101110010000", -- 11151 FREE #<CONS 0 11152>
 "00000000000000000010101110010001", -- 11152 FREE #<CONS 0 11153>
 "00000000000000000010101110010010", -- 11153 FREE #<CONS 0 11154>
 "00000000000000000010101110010011", -- 11154 FREE #<CONS 0 11155>
 "00000000000000000010101110010100", -- 11155 FREE #<CONS 0 11156>
 "00000000000000000010101110010101", -- 11156 FREE #<CONS 0 11157>
 "00000000000000000010101110010110", -- 11157 FREE #<CONS 0 11158>
 "00000000000000000010101110010111", -- 11158 FREE #<CONS 0 11159>
 "00000000000000000010101110011000", -- 11159 FREE #<CONS 0 11160>
 "00000000000000000010101110011001", -- 11160 FREE #<CONS 0 11161>
 "00000000000000000010101110011010", -- 11161 FREE #<CONS 0 11162>
 "00000000000000000010101110011011", -- 11162 FREE #<CONS 0 11163>
 "00000000000000000010101110011100", -- 11163 FREE #<CONS 0 11164>
 "00000000000000000010101110011101", -- 11164 FREE #<CONS 0 11165>
 "00000000000000000010101110011110", -- 11165 FREE #<CONS 0 11166>
 "00000000000000000010101110011111", -- 11166 FREE #<CONS 0 11167>
 "00000000000000000010101110100000", -- 11167 FREE #<CONS 0 11168>
 "00000000000000000010101110100001", -- 11168 FREE #<CONS 0 11169>
 "00000000000000000010101110100010", -- 11169 FREE #<CONS 0 11170>
 "00000000000000000010101110100011", -- 11170 FREE #<CONS 0 11171>
 "00000000000000000010101110100100", -- 11171 FREE #<CONS 0 11172>
 "00000000000000000010101110100101", -- 11172 FREE #<CONS 0 11173>
 "00000000000000000010101110100110", -- 11173 FREE #<CONS 0 11174>
 "00000000000000000010101110100111", -- 11174 FREE #<CONS 0 11175>
 "00000000000000000010101110101000", -- 11175 FREE #<CONS 0 11176>
 "00000000000000000010101110101001", -- 11176 FREE #<CONS 0 11177>
 "00000000000000000010101110101010", -- 11177 FREE #<CONS 0 11178>
 "00000000000000000010101110101011", -- 11178 FREE #<CONS 0 11179>
 "00000000000000000010101110101100", -- 11179 FREE #<CONS 0 11180>
 "00000000000000000010101110101101", -- 11180 FREE #<CONS 0 11181>
 "00000000000000000010101110101110", -- 11181 FREE #<CONS 0 11182>
 "00000000000000000010101110101111", -- 11182 FREE #<CONS 0 11183>
 "00000000000000000010101110110000", -- 11183 FREE #<CONS 0 11184>
 "00000000000000000010101110110001", -- 11184 FREE #<CONS 0 11185>
 "00000000000000000010101110110010", -- 11185 FREE #<CONS 0 11186>
 "00000000000000000010101110110011", -- 11186 FREE #<CONS 0 11187>
 "00000000000000000010101110110100", -- 11187 FREE #<CONS 0 11188>
 "00000000000000000010101110110101", -- 11188 FREE #<CONS 0 11189>
 "00000000000000000010101110110110", -- 11189 FREE #<CONS 0 11190>
 "00000000000000000010101110110111", -- 11190 FREE #<CONS 0 11191>
 "00000000000000000010101110111000", -- 11191 FREE #<CONS 0 11192>
 "00000000000000000010101110111001", -- 11192 FREE #<CONS 0 11193>
 "00000000000000000010101110111010", -- 11193 FREE #<CONS 0 11194>
 "00000000000000000010101110111011", -- 11194 FREE #<CONS 0 11195>
 "00000000000000000010101110111100", -- 11195 FREE #<CONS 0 11196>
 "00000000000000000010101110111101", -- 11196 FREE #<CONS 0 11197>
 "00000000000000000010101110111110", -- 11197 FREE #<CONS 0 11198>
 "00000000000000000010101110111111", -- 11198 FREE #<CONS 0 11199>
 "00000000000000000010101111000000", -- 11199 FREE #<CONS 0 11200>
 "00000000000000000010101111000001", -- 11200 FREE #<CONS 0 11201>
 "00000000000000000010101111000010", -- 11201 FREE #<CONS 0 11202>
 "00000000000000000010101111000011", -- 11202 FREE #<CONS 0 11203>
 "00000000000000000010101111000100", -- 11203 FREE #<CONS 0 11204>
 "00000000000000000010101111000101", -- 11204 FREE #<CONS 0 11205>
 "00000000000000000010101111000110", -- 11205 FREE #<CONS 0 11206>
 "00000000000000000010101111000111", -- 11206 FREE #<CONS 0 11207>
 "00000000000000000010101111001000", -- 11207 FREE #<CONS 0 11208>
 "00000000000000000010101111001001", -- 11208 FREE #<CONS 0 11209>
 "00000000000000000010101111001010", -- 11209 FREE #<CONS 0 11210>
 "00000000000000000010101111001011", -- 11210 FREE #<CONS 0 11211>
 "00000000000000000010101111001100", -- 11211 FREE #<CONS 0 11212>
 "00000000000000000010101111001101", -- 11212 FREE #<CONS 0 11213>
 "00000000000000000010101111001110", -- 11213 FREE #<CONS 0 11214>
 "00000000000000000010101111001111", -- 11214 FREE #<CONS 0 11215>
 "00000000000000000010101111010000", -- 11215 FREE #<CONS 0 11216>
 "00000000000000000010101111010001", -- 11216 FREE #<CONS 0 11217>
 "00000000000000000010101111010010", -- 11217 FREE #<CONS 0 11218>
 "00000000000000000010101111010011", -- 11218 FREE #<CONS 0 11219>
 "00000000000000000010101111010100", -- 11219 FREE #<CONS 0 11220>
 "00000000000000000010101111010101", -- 11220 FREE #<CONS 0 11221>
 "00000000000000000010101111010110", -- 11221 FREE #<CONS 0 11222>
 "00000000000000000010101111010111", -- 11222 FREE #<CONS 0 11223>
 "00000000000000000010101111011000", -- 11223 FREE #<CONS 0 11224>
 "00000000000000000010101111011001", -- 11224 FREE #<CONS 0 11225>
 "00000000000000000010101111011010", -- 11225 FREE #<CONS 0 11226>
 "00000000000000000010101111011011", -- 11226 FREE #<CONS 0 11227>
 "00000000000000000010101111011100", -- 11227 FREE #<CONS 0 11228>
 "00000000000000000010101111011101", -- 11228 FREE #<CONS 0 11229>
 "00000000000000000010101111011110", -- 11229 FREE #<CONS 0 11230>
 "00000000000000000010101111011111", -- 11230 FREE #<CONS 0 11231>
 "00000000000000000010101111100000", -- 11231 FREE #<CONS 0 11232>
 "00000000000000000010101111100001", -- 11232 FREE #<CONS 0 11233>
 "00000000000000000010101111100010", -- 11233 FREE #<CONS 0 11234>
 "00000000000000000010101111100011", -- 11234 FREE #<CONS 0 11235>
 "00000000000000000010101111100100", -- 11235 FREE #<CONS 0 11236>
 "00000000000000000010101111100101", -- 11236 FREE #<CONS 0 11237>
 "00000000000000000010101111100110", -- 11237 FREE #<CONS 0 11238>
 "00000000000000000010101111100111", -- 11238 FREE #<CONS 0 11239>
 "00000000000000000010101111101000", -- 11239 FREE #<CONS 0 11240>
 "00000000000000000010101111101001", -- 11240 FREE #<CONS 0 11241>
 "00000000000000000010101111101010", -- 11241 FREE #<CONS 0 11242>
 "00000000000000000010101111101011", -- 11242 FREE #<CONS 0 11243>
 "00000000000000000010101111101100", -- 11243 FREE #<CONS 0 11244>
 "00000000000000000010101111101101", -- 11244 FREE #<CONS 0 11245>
 "00000000000000000010101111101110", -- 11245 FREE #<CONS 0 11246>
 "00000000000000000010101111101111", -- 11246 FREE #<CONS 0 11247>
 "00000000000000000010101111110000", -- 11247 FREE #<CONS 0 11248>
 "00000000000000000010101111110001", -- 11248 FREE #<CONS 0 11249>
 "00000000000000000010101111110010", -- 11249 FREE #<CONS 0 11250>
 "00000000000000000010101111110011", -- 11250 FREE #<CONS 0 11251>
 "00000000000000000010101111110100", -- 11251 FREE #<CONS 0 11252>
 "00000000000000000010101111110101", -- 11252 FREE #<CONS 0 11253>
 "00000000000000000010101111110110", -- 11253 FREE #<CONS 0 11254>
 "00000000000000000010101111110111", -- 11254 FREE #<CONS 0 11255>
 "00000000000000000010101111111000", -- 11255 FREE #<CONS 0 11256>
 "00000000000000000010101111111001", -- 11256 FREE #<CONS 0 11257>
 "00000000000000000010101111111010", -- 11257 FREE #<CONS 0 11258>
 "00000000000000000010101111111011", -- 11258 FREE #<CONS 0 11259>
 "00000000000000000010101111111100", -- 11259 FREE #<CONS 0 11260>
 "00000000000000000010101111111101", -- 11260 FREE #<CONS 0 11261>
 "00000000000000000010101111111110", -- 11261 FREE #<CONS 0 11262>
 "00000000000000000010101111111111", -- 11262 FREE #<CONS 0 11263>
 "00000000000000000010110000000000", -- 11263 FREE #<CONS 0 11264>
 "00000000000000000010110000000001", -- 11264 FREE #<CONS 0 11265>
 "00000000000000000010110000000010", -- 11265 FREE #<CONS 0 11266>
 "00000000000000000010110000000011", -- 11266 FREE #<CONS 0 11267>
 "00000000000000000010110000000100", -- 11267 FREE #<CONS 0 11268>
 "00000000000000000010110000000101", -- 11268 FREE #<CONS 0 11269>
 "00000000000000000010110000000110", -- 11269 FREE #<CONS 0 11270>
 "00000000000000000010110000000111", -- 11270 FREE #<CONS 0 11271>
 "00000000000000000010110000001000", -- 11271 FREE #<CONS 0 11272>
 "00000000000000000010110000001001", -- 11272 FREE #<CONS 0 11273>
 "00000000000000000010110000001010", -- 11273 FREE #<CONS 0 11274>
 "00000000000000000010110000001011", -- 11274 FREE #<CONS 0 11275>
 "00000000000000000010110000001100", -- 11275 FREE #<CONS 0 11276>
 "00000000000000000010110000001101", -- 11276 FREE #<CONS 0 11277>
 "00000000000000000010110000001110", -- 11277 FREE #<CONS 0 11278>
 "00000000000000000010110000001111", -- 11278 FREE #<CONS 0 11279>
 "00000000000000000010110000010000", -- 11279 FREE #<CONS 0 11280>
 "00000000000000000010110000010001", -- 11280 FREE #<CONS 0 11281>
 "00000000000000000010110000010010", -- 11281 FREE #<CONS 0 11282>
 "00000000000000000010110000010011", -- 11282 FREE #<CONS 0 11283>
 "00000000000000000010110000010100", -- 11283 FREE #<CONS 0 11284>
 "00000000000000000010110000010101", -- 11284 FREE #<CONS 0 11285>
 "00000000000000000010110000010110", -- 11285 FREE #<CONS 0 11286>
 "00000000000000000010110000010111", -- 11286 FREE #<CONS 0 11287>
 "00000000000000000010110000011000", -- 11287 FREE #<CONS 0 11288>
 "00000000000000000010110000011001", -- 11288 FREE #<CONS 0 11289>
 "00000000000000000010110000011010", -- 11289 FREE #<CONS 0 11290>
 "00000000000000000010110000011011", -- 11290 FREE #<CONS 0 11291>
 "00000000000000000010110000011100", -- 11291 FREE #<CONS 0 11292>
 "00000000000000000010110000011101", -- 11292 FREE #<CONS 0 11293>
 "00000000000000000010110000011110", -- 11293 FREE #<CONS 0 11294>
 "00000000000000000010110000011111", -- 11294 FREE #<CONS 0 11295>
 "00000000000000000010110000100000", -- 11295 FREE #<CONS 0 11296>
 "00000000000000000010110000100001", -- 11296 FREE #<CONS 0 11297>
 "00000000000000000010110000100010", -- 11297 FREE #<CONS 0 11298>
 "00000000000000000010110000100011", -- 11298 FREE #<CONS 0 11299>
 "00000000000000000010110000100100", -- 11299 FREE #<CONS 0 11300>
 "00000000000000000010110000100101", -- 11300 FREE #<CONS 0 11301>
 "00000000000000000010110000100110", -- 11301 FREE #<CONS 0 11302>
 "00000000000000000010110000100111", -- 11302 FREE #<CONS 0 11303>
 "00000000000000000010110000101000", -- 11303 FREE #<CONS 0 11304>
 "00000000000000000010110000101001", -- 11304 FREE #<CONS 0 11305>
 "00000000000000000010110000101010", -- 11305 FREE #<CONS 0 11306>
 "00000000000000000010110000101011", -- 11306 FREE #<CONS 0 11307>
 "00000000000000000010110000101100", -- 11307 FREE #<CONS 0 11308>
 "00000000000000000010110000101101", -- 11308 FREE #<CONS 0 11309>
 "00000000000000000010110000101110", -- 11309 FREE #<CONS 0 11310>
 "00000000000000000010110000101111", -- 11310 FREE #<CONS 0 11311>
 "00000000000000000010110000110000", -- 11311 FREE #<CONS 0 11312>
 "00000000000000000010110000110001", -- 11312 FREE #<CONS 0 11313>
 "00000000000000000010110000110010", -- 11313 FREE #<CONS 0 11314>
 "00000000000000000010110000110011", -- 11314 FREE #<CONS 0 11315>
 "00000000000000000010110000110100", -- 11315 FREE #<CONS 0 11316>
 "00000000000000000010110000110101", -- 11316 FREE #<CONS 0 11317>
 "00000000000000000010110000110110", -- 11317 FREE #<CONS 0 11318>
 "00000000000000000010110000110111", -- 11318 FREE #<CONS 0 11319>
 "00000000000000000010110000111000", -- 11319 FREE #<CONS 0 11320>
 "00000000000000000010110000111001", -- 11320 FREE #<CONS 0 11321>
 "00000000000000000010110000111010", -- 11321 FREE #<CONS 0 11322>
 "00000000000000000010110000111011", -- 11322 FREE #<CONS 0 11323>
 "00000000000000000010110000111100", -- 11323 FREE #<CONS 0 11324>
 "00000000000000000010110000111101", -- 11324 FREE #<CONS 0 11325>
 "00000000000000000010110000111110", -- 11325 FREE #<CONS 0 11326>
 "00000000000000000010110000111111", -- 11326 FREE #<CONS 0 11327>
 "00000000000000000010110001000000", -- 11327 FREE #<CONS 0 11328>
 "00000000000000000010110001000001", -- 11328 FREE #<CONS 0 11329>
 "00000000000000000010110001000010", -- 11329 FREE #<CONS 0 11330>
 "00000000000000000010110001000011", -- 11330 FREE #<CONS 0 11331>
 "00000000000000000010110001000100", -- 11331 FREE #<CONS 0 11332>
 "00000000000000000010110001000101", -- 11332 FREE #<CONS 0 11333>
 "00000000000000000010110001000110", -- 11333 FREE #<CONS 0 11334>
 "00000000000000000010110001000111", -- 11334 FREE #<CONS 0 11335>
 "00000000000000000010110001001000", -- 11335 FREE #<CONS 0 11336>
 "00000000000000000010110001001001", -- 11336 FREE #<CONS 0 11337>
 "00000000000000000010110001001010", -- 11337 FREE #<CONS 0 11338>
 "00000000000000000010110001001011", -- 11338 FREE #<CONS 0 11339>
 "00000000000000000010110001001100", -- 11339 FREE #<CONS 0 11340>
 "00000000000000000010110001001101", -- 11340 FREE #<CONS 0 11341>
 "00000000000000000010110001001110", -- 11341 FREE #<CONS 0 11342>
 "00000000000000000010110001001111", -- 11342 FREE #<CONS 0 11343>
 "00000000000000000010110001010000", -- 11343 FREE #<CONS 0 11344>
 "00000000000000000010110001010001", -- 11344 FREE #<CONS 0 11345>
 "00000000000000000010110001010010", -- 11345 FREE #<CONS 0 11346>
 "00000000000000000010110001010011", -- 11346 FREE #<CONS 0 11347>
 "00000000000000000010110001010100", -- 11347 FREE #<CONS 0 11348>
 "00000000000000000010110001010101", -- 11348 FREE #<CONS 0 11349>
 "00000000000000000010110001010110", -- 11349 FREE #<CONS 0 11350>
 "00000000000000000010110001010111", -- 11350 FREE #<CONS 0 11351>
 "00000000000000000010110001011000", -- 11351 FREE #<CONS 0 11352>
 "00000000000000000010110001011001", -- 11352 FREE #<CONS 0 11353>
 "00000000000000000010110001011010", -- 11353 FREE #<CONS 0 11354>
 "00000000000000000010110001011011", -- 11354 FREE #<CONS 0 11355>
 "00000000000000000010110001011100", -- 11355 FREE #<CONS 0 11356>
 "00000000000000000010110001011101", -- 11356 FREE #<CONS 0 11357>
 "00000000000000000010110001011110", -- 11357 FREE #<CONS 0 11358>
 "00000000000000000010110001011111", -- 11358 FREE #<CONS 0 11359>
 "00000000000000000010110001100000", -- 11359 FREE #<CONS 0 11360>
 "00000000000000000010110001100001", -- 11360 FREE #<CONS 0 11361>
 "00000000000000000010110001100010", -- 11361 FREE #<CONS 0 11362>
 "00000000000000000010110001100011", -- 11362 FREE #<CONS 0 11363>
 "00000000000000000010110001100100", -- 11363 FREE #<CONS 0 11364>
 "00000000000000000010110001100101", -- 11364 FREE #<CONS 0 11365>
 "00000000000000000010110001100110", -- 11365 FREE #<CONS 0 11366>
 "00000000000000000010110001100111", -- 11366 FREE #<CONS 0 11367>
 "00000000000000000010110001101000", -- 11367 FREE #<CONS 0 11368>
 "00000000000000000010110001101001", -- 11368 FREE #<CONS 0 11369>
 "00000000000000000010110001101010", -- 11369 FREE #<CONS 0 11370>
 "00000000000000000010110001101011", -- 11370 FREE #<CONS 0 11371>
 "00000000000000000010110001101100", -- 11371 FREE #<CONS 0 11372>
 "00000000000000000010110001101101", -- 11372 FREE #<CONS 0 11373>
 "00000000000000000010110001101110", -- 11373 FREE #<CONS 0 11374>
 "00000000000000000010110001101111", -- 11374 FREE #<CONS 0 11375>
 "00000000000000000010110001110000", -- 11375 FREE #<CONS 0 11376>
 "00000000000000000010110001110001", -- 11376 FREE #<CONS 0 11377>
 "00000000000000000010110001110010", -- 11377 FREE #<CONS 0 11378>
 "00000000000000000010110001110011", -- 11378 FREE #<CONS 0 11379>
 "00000000000000000010110001110100", -- 11379 FREE #<CONS 0 11380>
 "00000000000000000010110001110101", -- 11380 FREE #<CONS 0 11381>
 "00000000000000000010110001110110", -- 11381 FREE #<CONS 0 11382>
 "00000000000000000010110001110111", -- 11382 FREE #<CONS 0 11383>
 "00000000000000000010110001111000", -- 11383 FREE #<CONS 0 11384>
 "00000000000000000010110001111001", -- 11384 FREE #<CONS 0 11385>
 "00000000000000000010110001111010", -- 11385 FREE #<CONS 0 11386>
 "00000000000000000010110001111011", -- 11386 FREE #<CONS 0 11387>
 "00000000000000000010110001111100", -- 11387 FREE #<CONS 0 11388>
 "00000000000000000010110001111101", -- 11388 FREE #<CONS 0 11389>
 "00000000000000000010110001111110", -- 11389 FREE #<CONS 0 11390>
 "00000000000000000010110001111111", -- 11390 FREE #<CONS 0 11391>
 "00000000000000000010110010000000", -- 11391 FREE #<CONS 0 11392>
 "00000000000000000010110010000001", -- 11392 FREE #<CONS 0 11393>
 "00000000000000000010110010000010", -- 11393 FREE #<CONS 0 11394>
 "00000000000000000010110010000011", -- 11394 FREE #<CONS 0 11395>
 "00000000000000000010110010000100", -- 11395 FREE #<CONS 0 11396>
 "00000000000000000010110010000101", -- 11396 FREE #<CONS 0 11397>
 "00000000000000000010110010000110", -- 11397 FREE #<CONS 0 11398>
 "00000000000000000010110010000111", -- 11398 FREE #<CONS 0 11399>
 "00000000000000000010110010001000", -- 11399 FREE #<CONS 0 11400>
 "00000000000000000010110010001001", -- 11400 FREE #<CONS 0 11401>
 "00000000000000000010110010001010", -- 11401 FREE #<CONS 0 11402>
 "00000000000000000010110010001011", -- 11402 FREE #<CONS 0 11403>
 "00000000000000000010110010001100", -- 11403 FREE #<CONS 0 11404>
 "00000000000000000010110010001101", -- 11404 FREE #<CONS 0 11405>
 "00000000000000000010110010001110", -- 11405 FREE #<CONS 0 11406>
 "00000000000000000010110010001111", -- 11406 FREE #<CONS 0 11407>
 "00000000000000000010110010010000", -- 11407 FREE #<CONS 0 11408>
 "00000000000000000010110010010001", -- 11408 FREE #<CONS 0 11409>
 "00000000000000000010110010010010", -- 11409 FREE #<CONS 0 11410>
 "00000000000000000010110010010011", -- 11410 FREE #<CONS 0 11411>
 "00000000000000000010110010010100", -- 11411 FREE #<CONS 0 11412>
 "00000000000000000010110010010101", -- 11412 FREE #<CONS 0 11413>
 "00000000000000000010110010010110", -- 11413 FREE #<CONS 0 11414>
 "00000000000000000010110010010111", -- 11414 FREE #<CONS 0 11415>
 "00000000000000000010110010011000", -- 11415 FREE #<CONS 0 11416>
 "00000000000000000010110010011001", -- 11416 FREE #<CONS 0 11417>
 "00000000000000000010110010011010", -- 11417 FREE #<CONS 0 11418>
 "00000000000000000010110010011011", -- 11418 FREE #<CONS 0 11419>
 "00000000000000000010110010011100", -- 11419 FREE #<CONS 0 11420>
 "00000000000000000010110010011101", -- 11420 FREE #<CONS 0 11421>
 "00000000000000000010110010011110", -- 11421 FREE #<CONS 0 11422>
 "00000000000000000010110010011111", -- 11422 FREE #<CONS 0 11423>
 "00000000000000000010110010100000", -- 11423 FREE #<CONS 0 11424>
 "00000000000000000010110010100001", -- 11424 FREE #<CONS 0 11425>
 "00000000000000000010110010100010", -- 11425 FREE #<CONS 0 11426>
 "00000000000000000010110010100011", -- 11426 FREE #<CONS 0 11427>
 "00000000000000000010110010100100", -- 11427 FREE #<CONS 0 11428>
 "00000000000000000010110010100101", -- 11428 FREE #<CONS 0 11429>
 "00000000000000000010110010100110", -- 11429 FREE #<CONS 0 11430>
 "00000000000000000010110010100111", -- 11430 FREE #<CONS 0 11431>
 "00000000000000000010110010101000", -- 11431 FREE #<CONS 0 11432>
 "00000000000000000010110010101001", -- 11432 FREE #<CONS 0 11433>
 "00000000000000000010110010101010", -- 11433 FREE #<CONS 0 11434>
 "00000000000000000010110010101011", -- 11434 FREE #<CONS 0 11435>
 "00000000000000000010110010101100", -- 11435 FREE #<CONS 0 11436>
 "00000000000000000010110010101101", -- 11436 FREE #<CONS 0 11437>
 "00000000000000000010110010101110", -- 11437 FREE #<CONS 0 11438>
 "00000000000000000010110010101111", -- 11438 FREE #<CONS 0 11439>
 "00000000000000000010110010110000", -- 11439 FREE #<CONS 0 11440>
 "00000000000000000010110010110001", -- 11440 FREE #<CONS 0 11441>
 "00000000000000000010110010110010", -- 11441 FREE #<CONS 0 11442>
 "00000000000000000010110010110011", -- 11442 FREE #<CONS 0 11443>
 "00000000000000000010110010110100", -- 11443 FREE #<CONS 0 11444>
 "00000000000000000010110010110101", -- 11444 FREE #<CONS 0 11445>
 "00000000000000000010110010110110", -- 11445 FREE #<CONS 0 11446>
 "00000000000000000010110010110111", -- 11446 FREE #<CONS 0 11447>
 "00000000000000000010110010111000", -- 11447 FREE #<CONS 0 11448>
 "00000000000000000010110010111001", -- 11448 FREE #<CONS 0 11449>
 "00000000000000000010110010111010", -- 11449 FREE #<CONS 0 11450>
 "00000000000000000010110010111011", -- 11450 FREE #<CONS 0 11451>
 "00000000000000000010110010111100", -- 11451 FREE #<CONS 0 11452>
 "00000000000000000010110010111101", -- 11452 FREE #<CONS 0 11453>
 "00000000000000000010110010111110", -- 11453 FREE #<CONS 0 11454>
 "00000000000000000010110010111111", -- 11454 FREE #<CONS 0 11455>
 "00000000000000000010110011000000", -- 11455 FREE #<CONS 0 11456>
 "00000000000000000010110011000001", -- 11456 FREE #<CONS 0 11457>
 "00000000000000000010110011000010", -- 11457 FREE #<CONS 0 11458>
 "00000000000000000010110011000011", -- 11458 FREE #<CONS 0 11459>
 "00000000000000000010110011000100", -- 11459 FREE #<CONS 0 11460>
 "00000000000000000010110011000101", -- 11460 FREE #<CONS 0 11461>
 "00000000000000000010110011000110", -- 11461 FREE #<CONS 0 11462>
 "00000000000000000010110011000111", -- 11462 FREE #<CONS 0 11463>
 "00000000000000000010110011001000", -- 11463 FREE #<CONS 0 11464>
 "00000000000000000010110011001001", -- 11464 FREE #<CONS 0 11465>
 "00000000000000000010110011001010", -- 11465 FREE #<CONS 0 11466>
 "00000000000000000010110011001011", -- 11466 FREE #<CONS 0 11467>
 "00000000000000000010110011001100", -- 11467 FREE #<CONS 0 11468>
 "00000000000000000010110011001101", -- 11468 FREE #<CONS 0 11469>
 "00000000000000000010110011001110", -- 11469 FREE #<CONS 0 11470>
 "00000000000000000010110011001111", -- 11470 FREE #<CONS 0 11471>
 "00000000000000000010110011010000", -- 11471 FREE #<CONS 0 11472>
 "00000000000000000010110011010001", -- 11472 FREE #<CONS 0 11473>
 "00000000000000000010110011010010", -- 11473 FREE #<CONS 0 11474>
 "00000000000000000010110011010011", -- 11474 FREE #<CONS 0 11475>
 "00000000000000000010110011010100", -- 11475 FREE #<CONS 0 11476>
 "00000000000000000010110011010101", -- 11476 FREE #<CONS 0 11477>
 "00000000000000000010110011010110", -- 11477 FREE #<CONS 0 11478>
 "00000000000000000010110011010111", -- 11478 FREE #<CONS 0 11479>
 "00000000000000000010110011011000", -- 11479 FREE #<CONS 0 11480>
 "00000000000000000010110011011001", -- 11480 FREE #<CONS 0 11481>
 "00000000000000000010110011011010", -- 11481 FREE #<CONS 0 11482>
 "00000000000000000010110011011011", -- 11482 FREE #<CONS 0 11483>
 "00000000000000000010110011011100", -- 11483 FREE #<CONS 0 11484>
 "00000000000000000010110011011101", -- 11484 FREE #<CONS 0 11485>
 "00000000000000000010110011011110", -- 11485 FREE #<CONS 0 11486>
 "00000000000000000010110011011111", -- 11486 FREE #<CONS 0 11487>
 "00000000000000000010110011100000", -- 11487 FREE #<CONS 0 11488>
 "00000000000000000010110011100001", -- 11488 FREE #<CONS 0 11489>
 "00000000000000000010110011100010", -- 11489 FREE #<CONS 0 11490>
 "00000000000000000010110011100011", -- 11490 FREE #<CONS 0 11491>
 "00000000000000000010110011100100", -- 11491 FREE #<CONS 0 11492>
 "00000000000000000010110011100101", -- 11492 FREE #<CONS 0 11493>
 "00000000000000000010110011100110", -- 11493 FREE #<CONS 0 11494>
 "00000000000000000010110011100111", -- 11494 FREE #<CONS 0 11495>
 "00000000000000000010110011101000", -- 11495 FREE #<CONS 0 11496>
 "00000000000000000010110011101001", -- 11496 FREE #<CONS 0 11497>
 "00000000000000000010110011101010", -- 11497 FREE #<CONS 0 11498>
 "00000000000000000010110011101011", -- 11498 FREE #<CONS 0 11499>
 "00000000000000000010110011101100", -- 11499 FREE #<CONS 0 11500>
 "00000000000000000010110011101101", -- 11500 FREE #<CONS 0 11501>
 "00000000000000000010110011101110", -- 11501 FREE #<CONS 0 11502>
 "00000000000000000010110011101111", -- 11502 FREE #<CONS 0 11503>
 "00000000000000000010110011110000", -- 11503 FREE #<CONS 0 11504>
 "00000000000000000010110011110001", -- 11504 FREE #<CONS 0 11505>
 "00000000000000000010110011110010", -- 11505 FREE #<CONS 0 11506>
 "00000000000000000010110011110011", -- 11506 FREE #<CONS 0 11507>
 "00000000000000000010110011110100", -- 11507 FREE #<CONS 0 11508>
 "00000000000000000010110011110101", -- 11508 FREE #<CONS 0 11509>
 "00000000000000000010110011110110", -- 11509 FREE #<CONS 0 11510>
 "00000000000000000010110011110111", -- 11510 FREE #<CONS 0 11511>
 "00000000000000000010110011111000", -- 11511 FREE #<CONS 0 11512>
 "00000000000000000010110011111001", -- 11512 FREE #<CONS 0 11513>
 "00000000000000000010110011111010", -- 11513 FREE #<CONS 0 11514>
 "00000000000000000010110011111011", -- 11514 FREE #<CONS 0 11515>
 "00000000000000000010110011111100", -- 11515 FREE #<CONS 0 11516>
 "00000000000000000010110011111101", -- 11516 FREE #<CONS 0 11517>
 "00000000000000000010110011111110", -- 11517 FREE #<CONS 0 11518>
 "00000000000000000010110011111111", -- 11518 FREE #<CONS 0 11519>
 "00000000000000000010110100000000", -- 11519 FREE #<CONS 0 11520>
 "00000000000000000010110100000001", -- 11520 FREE #<CONS 0 11521>
 "00000000000000000010110100000010", -- 11521 FREE #<CONS 0 11522>
 "00000000000000000010110100000011", -- 11522 FREE #<CONS 0 11523>
 "00000000000000000010110100000100", -- 11523 FREE #<CONS 0 11524>
 "00000000000000000010110100000101", -- 11524 FREE #<CONS 0 11525>
 "00000000000000000010110100000110", -- 11525 FREE #<CONS 0 11526>
 "00000000000000000010110100000111", -- 11526 FREE #<CONS 0 11527>
 "00000000000000000010110100001000", -- 11527 FREE #<CONS 0 11528>
 "00000000000000000010110100001001", -- 11528 FREE #<CONS 0 11529>
 "00000000000000000010110100001010", -- 11529 FREE #<CONS 0 11530>
 "00000000000000000010110100001011", -- 11530 FREE #<CONS 0 11531>
 "00000000000000000010110100001100", -- 11531 FREE #<CONS 0 11532>
 "00000000000000000010110100001101", -- 11532 FREE #<CONS 0 11533>
 "00000000000000000010110100001110", -- 11533 FREE #<CONS 0 11534>
 "00000000000000000010110100001111", -- 11534 FREE #<CONS 0 11535>
 "00000000000000000010110100010000", -- 11535 FREE #<CONS 0 11536>
 "00000000000000000010110100010001", -- 11536 FREE #<CONS 0 11537>
 "00000000000000000010110100010010", -- 11537 FREE #<CONS 0 11538>
 "00000000000000000010110100010011", -- 11538 FREE #<CONS 0 11539>
 "00000000000000000010110100010100", -- 11539 FREE #<CONS 0 11540>
 "00000000000000000010110100010101", -- 11540 FREE #<CONS 0 11541>
 "00000000000000000010110100010110", -- 11541 FREE #<CONS 0 11542>
 "00000000000000000010110100010111", -- 11542 FREE #<CONS 0 11543>
 "00000000000000000010110100011000", -- 11543 FREE #<CONS 0 11544>
 "00000000000000000010110100011001", -- 11544 FREE #<CONS 0 11545>
 "00000000000000000010110100011010", -- 11545 FREE #<CONS 0 11546>
 "00000000000000000010110100011011", -- 11546 FREE #<CONS 0 11547>
 "00000000000000000010110100011100", -- 11547 FREE #<CONS 0 11548>
 "00000000000000000010110100011101", -- 11548 FREE #<CONS 0 11549>
 "00000000000000000010110100011110", -- 11549 FREE #<CONS 0 11550>
 "00000000000000000010110100011111", -- 11550 FREE #<CONS 0 11551>
 "00000000000000000010110100100000", -- 11551 FREE #<CONS 0 11552>
 "00000000000000000010110100100001", -- 11552 FREE #<CONS 0 11553>
 "00000000000000000010110100100010", -- 11553 FREE #<CONS 0 11554>
 "00000000000000000010110100100011", -- 11554 FREE #<CONS 0 11555>
 "00000000000000000010110100100100", -- 11555 FREE #<CONS 0 11556>
 "00000000000000000010110100100101", -- 11556 FREE #<CONS 0 11557>
 "00000000000000000010110100100110", -- 11557 FREE #<CONS 0 11558>
 "00000000000000000010110100100111", -- 11558 FREE #<CONS 0 11559>
 "00000000000000000010110100101000", -- 11559 FREE #<CONS 0 11560>
 "00000000000000000010110100101001", -- 11560 FREE #<CONS 0 11561>
 "00000000000000000010110100101010", -- 11561 FREE #<CONS 0 11562>
 "00000000000000000010110100101011", -- 11562 FREE #<CONS 0 11563>
 "00000000000000000010110100101100", -- 11563 FREE #<CONS 0 11564>
 "00000000000000000010110100101101", -- 11564 FREE #<CONS 0 11565>
 "00000000000000000010110100101110", -- 11565 FREE #<CONS 0 11566>
 "00000000000000000010110100101111", -- 11566 FREE #<CONS 0 11567>
 "00000000000000000010110100110000", -- 11567 FREE #<CONS 0 11568>
 "00000000000000000010110100110001", -- 11568 FREE #<CONS 0 11569>
 "00000000000000000010110100110010", -- 11569 FREE #<CONS 0 11570>
 "00000000000000000010110100110011", -- 11570 FREE #<CONS 0 11571>
 "00000000000000000010110100110100", -- 11571 FREE #<CONS 0 11572>
 "00000000000000000010110100110101", -- 11572 FREE #<CONS 0 11573>
 "00000000000000000010110100110110", -- 11573 FREE #<CONS 0 11574>
 "00000000000000000010110100110111", -- 11574 FREE #<CONS 0 11575>
 "00000000000000000010110100111000", -- 11575 FREE #<CONS 0 11576>
 "00000000000000000010110100111001", -- 11576 FREE #<CONS 0 11577>
 "00000000000000000010110100111010", -- 11577 FREE #<CONS 0 11578>
 "00000000000000000010110100111011", -- 11578 FREE #<CONS 0 11579>
 "00000000000000000010110100111100", -- 11579 FREE #<CONS 0 11580>
 "00000000000000000010110100111101", -- 11580 FREE #<CONS 0 11581>
 "00000000000000000010110100111110", -- 11581 FREE #<CONS 0 11582>
 "00000000000000000010110100111111", -- 11582 FREE #<CONS 0 11583>
 "00000000000000000010110101000000", -- 11583 FREE #<CONS 0 11584>
 "00000000000000000010110101000001", -- 11584 FREE #<CONS 0 11585>
 "00000000000000000010110101000010", -- 11585 FREE #<CONS 0 11586>
 "00000000000000000010110101000011", -- 11586 FREE #<CONS 0 11587>
 "00000000000000000010110101000100", -- 11587 FREE #<CONS 0 11588>
 "00000000000000000010110101000101", -- 11588 FREE #<CONS 0 11589>
 "00000000000000000010110101000110", -- 11589 FREE #<CONS 0 11590>
 "00000000000000000010110101000111", -- 11590 FREE #<CONS 0 11591>
 "00000000000000000010110101001000", -- 11591 FREE #<CONS 0 11592>
 "00000000000000000010110101001001", -- 11592 FREE #<CONS 0 11593>
 "00000000000000000010110101001010", -- 11593 FREE #<CONS 0 11594>
 "00000000000000000010110101001011", -- 11594 FREE #<CONS 0 11595>
 "00000000000000000010110101001100", -- 11595 FREE #<CONS 0 11596>
 "00000000000000000010110101001101", -- 11596 FREE #<CONS 0 11597>
 "00000000000000000010110101001110", -- 11597 FREE #<CONS 0 11598>
 "00000000000000000010110101001111", -- 11598 FREE #<CONS 0 11599>
 "00000000000000000010110101010000", -- 11599 FREE #<CONS 0 11600>
 "00000000000000000010110101010001", -- 11600 FREE #<CONS 0 11601>
 "00000000000000000010110101010010", -- 11601 FREE #<CONS 0 11602>
 "00000000000000000010110101010011", -- 11602 FREE #<CONS 0 11603>
 "00000000000000000010110101010100", -- 11603 FREE #<CONS 0 11604>
 "00000000000000000010110101010101", -- 11604 FREE #<CONS 0 11605>
 "00000000000000000010110101010110", -- 11605 FREE #<CONS 0 11606>
 "00000000000000000010110101010111", -- 11606 FREE #<CONS 0 11607>
 "00000000000000000010110101011000", -- 11607 FREE #<CONS 0 11608>
 "00000000000000000010110101011001", -- 11608 FREE #<CONS 0 11609>
 "00000000000000000010110101011010", -- 11609 FREE #<CONS 0 11610>
 "00000000000000000010110101011011", -- 11610 FREE #<CONS 0 11611>
 "00000000000000000010110101011100", -- 11611 FREE #<CONS 0 11612>
 "00000000000000000010110101011101", -- 11612 FREE #<CONS 0 11613>
 "00000000000000000010110101011110", -- 11613 FREE #<CONS 0 11614>
 "00000000000000000010110101011111", -- 11614 FREE #<CONS 0 11615>
 "00000000000000000010110101100000", -- 11615 FREE #<CONS 0 11616>
 "00000000000000000010110101100001", -- 11616 FREE #<CONS 0 11617>
 "00000000000000000010110101100010", -- 11617 FREE #<CONS 0 11618>
 "00000000000000000010110101100011", -- 11618 FREE #<CONS 0 11619>
 "00000000000000000010110101100100", -- 11619 FREE #<CONS 0 11620>
 "00000000000000000010110101100101", -- 11620 FREE #<CONS 0 11621>
 "00000000000000000010110101100110", -- 11621 FREE #<CONS 0 11622>
 "00000000000000000010110101100111", -- 11622 FREE #<CONS 0 11623>
 "00000000000000000010110101101000", -- 11623 FREE #<CONS 0 11624>
 "00000000000000000010110101101001", -- 11624 FREE #<CONS 0 11625>
 "00000000000000000010110101101010", -- 11625 FREE #<CONS 0 11626>
 "00000000000000000010110101101011", -- 11626 FREE #<CONS 0 11627>
 "00000000000000000010110101101100", -- 11627 FREE #<CONS 0 11628>
 "00000000000000000010110101101101", -- 11628 FREE #<CONS 0 11629>
 "00000000000000000010110101101110", -- 11629 FREE #<CONS 0 11630>
 "00000000000000000010110101101111", -- 11630 FREE #<CONS 0 11631>
 "00000000000000000010110101110000", -- 11631 FREE #<CONS 0 11632>
 "00000000000000000010110101110001", -- 11632 FREE #<CONS 0 11633>
 "00000000000000000010110101110010", -- 11633 FREE #<CONS 0 11634>
 "00000000000000000010110101110011", -- 11634 FREE #<CONS 0 11635>
 "00000000000000000010110101110100", -- 11635 FREE #<CONS 0 11636>
 "00000000000000000010110101110101", -- 11636 FREE #<CONS 0 11637>
 "00000000000000000010110101110110", -- 11637 FREE #<CONS 0 11638>
 "00000000000000000010110101110111", -- 11638 FREE #<CONS 0 11639>
 "00000000000000000010110101111000", -- 11639 FREE #<CONS 0 11640>
 "00000000000000000010110101111001", -- 11640 FREE #<CONS 0 11641>
 "00000000000000000010110101111010", -- 11641 FREE #<CONS 0 11642>
 "00000000000000000010110101111011", -- 11642 FREE #<CONS 0 11643>
 "00000000000000000010110101111100", -- 11643 FREE #<CONS 0 11644>
 "00000000000000000010110101111101", -- 11644 FREE #<CONS 0 11645>
 "00000000000000000010110101111110", -- 11645 FREE #<CONS 0 11646>
 "00000000000000000010110101111111", -- 11646 FREE #<CONS 0 11647>
 "00000000000000000010110110000000", -- 11647 FREE #<CONS 0 11648>
 "00000000000000000010110110000001", -- 11648 FREE #<CONS 0 11649>
 "00000000000000000010110110000010", -- 11649 FREE #<CONS 0 11650>
 "00000000000000000010110110000011", -- 11650 FREE #<CONS 0 11651>
 "00000000000000000010110110000100", -- 11651 FREE #<CONS 0 11652>
 "00000000000000000010110110000101", -- 11652 FREE #<CONS 0 11653>
 "00000000000000000010110110000110", -- 11653 FREE #<CONS 0 11654>
 "00000000000000000010110110000111", -- 11654 FREE #<CONS 0 11655>
 "00000000000000000010110110001000", -- 11655 FREE #<CONS 0 11656>
 "00000000000000000010110110001001", -- 11656 FREE #<CONS 0 11657>
 "00000000000000000010110110001010", -- 11657 FREE #<CONS 0 11658>
 "00000000000000000010110110001011", -- 11658 FREE #<CONS 0 11659>
 "00000000000000000010110110001100", -- 11659 FREE #<CONS 0 11660>
 "00000000000000000010110110001101", -- 11660 FREE #<CONS 0 11661>
 "00000000000000000010110110001110", -- 11661 FREE #<CONS 0 11662>
 "00000000000000000010110110001111", -- 11662 FREE #<CONS 0 11663>
 "00000000000000000010110110010000", -- 11663 FREE #<CONS 0 11664>
 "00000000000000000010110110010001", -- 11664 FREE #<CONS 0 11665>
 "00000000000000000010110110010010", -- 11665 FREE #<CONS 0 11666>
 "00000000000000000010110110010011", -- 11666 FREE #<CONS 0 11667>
 "00000000000000000010110110010100", -- 11667 FREE #<CONS 0 11668>
 "00000000000000000010110110010101", -- 11668 FREE #<CONS 0 11669>
 "00000000000000000010110110010110", -- 11669 FREE #<CONS 0 11670>
 "00000000000000000010110110010111", -- 11670 FREE #<CONS 0 11671>
 "00000000000000000010110110011000", -- 11671 FREE #<CONS 0 11672>
 "00000000000000000010110110011001", -- 11672 FREE #<CONS 0 11673>
 "00000000000000000010110110011010", -- 11673 FREE #<CONS 0 11674>
 "00000000000000000010110110011011", -- 11674 FREE #<CONS 0 11675>
 "00000000000000000010110110011100", -- 11675 FREE #<CONS 0 11676>
 "00000000000000000010110110011101", -- 11676 FREE #<CONS 0 11677>
 "00000000000000000010110110011110", -- 11677 FREE #<CONS 0 11678>
 "00000000000000000010110110011111", -- 11678 FREE #<CONS 0 11679>
 "00000000000000000010110110100000", -- 11679 FREE #<CONS 0 11680>
 "00000000000000000010110110100001", -- 11680 FREE #<CONS 0 11681>
 "00000000000000000010110110100010", -- 11681 FREE #<CONS 0 11682>
 "00000000000000000010110110100011", -- 11682 FREE #<CONS 0 11683>
 "00000000000000000010110110100100", -- 11683 FREE #<CONS 0 11684>
 "00000000000000000010110110100101", -- 11684 FREE #<CONS 0 11685>
 "00000000000000000010110110100110", -- 11685 FREE #<CONS 0 11686>
 "00000000000000000010110110100111", -- 11686 FREE #<CONS 0 11687>
 "00000000000000000010110110101000", -- 11687 FREE #<CONS 0 11688>
 "00000000000000000010110110101001", -- 11688 FREE #<CONS 0 11689>
 "00000000000000000010110110101010", -- 11689 FREE #<CONS 0 11690>
 "00000000000000000010110110101011", -- 11690 FREE #<CONS 0 11691>
 "00000000000000000010110110101100", -- 11691 FREE #<CONS 0 11692>
 "00000000000000000010110110101101", -- 11692 FREE #<CONS 0 11693>
 "00000000000000000010110110101110", -- 11693 FREE #<CONS 0 11694>
 "00000000000000000010110110101111", -- 11694 FREE #<CONS 0 11695>
 "00000000000000000010110110110000", -- 11695 FREE #<CONS 0 11696>
 "00000000000000000010110110110001", -- 11696 FREE #<CONS 0 11697>
 "00000000000000000010110110110010", -- 11697 FREE #<CONS 0 11698>
 "00000000000000000010110110110011", -- 11698 FREE #<CONS 0 11699>
 "00000000000000000010110110110100", -- 11699 FREE #<CONS 0 11700>
 "00000000000000000010110110110101", -- 11700 FREE #<CONS 0 11701>
 "00000000000000000010110110110110", -- 11701 FREE #<CONS 0 11702>
 "00000000000000000010110110110111", -- 11702 FREE #<CONS 0 11703>
 "00000000000000000010110110111000", -- 11703 FREE #<CONS 0 11704>
 "00000000000000000010110110111001", -- 11704 FREE #<CONS 0 11705>
 "00000000000000000010110110111010", -- 11705 FREE #<CONS 0 11706>
 "00000000000000000010110110111011", -- 11706 FREE #<CONS 0 11707>
 "00000000000000000010110110111100", -- 11707 FREE #<CONS 0 11708>
 "00000000000000000010110110111101", -- 11708 FREE #<CONS 0 11709>
 "00000000000000000010110110111110", -- 11709 FREE #<CONS 0 11710>
 "00000000000000000010110110111111", -- 11710 FREE #<CONS 0 11711>
 "00000000000000000010110111000000", -- 11711 FREE #<CONS 0 11712>
 "00000000000000000010110111000001", -- 11712 FREE #<CONS 0 11713>
 "00000000000000000010110111000010", -- 11713 FREE #<CONS 0 11714>
 "00000000000000000010110111000011", -- 11714 FREE #<CONS 0 11715>
 "00000000000000000010110111000100", -- 11715 FREE #<CONS 0 11716>
 "00000000000000000010110111000101", -- 11716 FREE #<CONS 0 11717>
 "00000000000000000010110111000110", -- 11717 FREE #<CONS 0 11718>
 "00000000000000000010110111000111", -- 11718 FREE #<CONS 0 11719>
 "00000000000000000010110111001000", -- 11719 FREE #<CONS 0 11720>
 "00000000000000000010110111001001", -- 11720 FREE #<CONS 0 11721>
 "00000000000000000010110111001010", -- 11721 FREE #<CONS 0 11722>
 "00000000000000000010110111001011", -- 11722 FREE #<CONS 0 11723>
 "00000000000000000010110111001100", -- 11723 FREE #<CONS 0 11724>
 "00000000000000000010110111001101", -- 11724 FREE #<CONS 0 11725>
 "00000000000000000010110111001110", -- 11725 FREE #<CONS 0 11726>
 "00000000000000000010110111001111", -- 11726 FREE #<CONS 0 11727>
 "00000000000000000010110111010000", -- 11727 FREE #<CONS 0 11728>
 "00000000000000000010110111010001", -- 11728 FREE #<CONS 0 11729>
 "00000000000000000010110111010010", -- 11729 FREE #<CONS 0 11730>
 "00000000000000000010110111010011", -- 11730 FREE #<CONS 0 11731>
 "00000000000000000010110111010100", -- 11731 FREE #<CONS 0 11732>
 "00000000000000000010110111010101", -- 11732 FREE #<CONS 0 11733>
 "00000000000000000010110111010110", -- 11733 FREE #<CONS 0 11734>
 "00000000000000000010110111010111", -- 11734 FREE #<CONS 0 11735>
 "00000000000000000010110111011000", -- 11735 FREE #<CONS 0 11736>
 "00000000000000000010110111011001", -- 11736 FREE #<CONS 0 11737>
 "00000000000000000010110111011010", -- 11737 FREE #<CONS 0 11738>
 "00000000000000000010110111011011", -- 11738 FREE #<CONS 0 11739>
 "00000000000000000010110111011100", -- 11739 FREE #<CONS 0 11740>
 "00000000000000000010110111011101", -- 11740 FREE #<CONS 0 11741>
 "00000000000000000010110111011110", -- 11741 FREE #<CONS 0 11742>
 "00000000000000000010110111011111", -- 11742 FREE #<CONS 0 11743>
 "00000000000000000010110111100000", -- 11743 FREE #<CONS 0 11744>
 "00000000000000000010110111100001", -- 11744 FREE #<CONS 0 11745>
 "00000000000000000010110111100010", -- 11745 FREE #<CONS 0 11746>
 "00000000000000000010110111100011", -- 11746 FREE #<CONS 0 11747>
 "00000000000000000010110111100100", -- 11747 FREE #<CONS 0 11748>
 "00000000000000000010110111100101", -- 11748 FREE #<CONS 0 11749>
 "00000000000000000010110111100110", -- 11749 FREE #<CONS 0 11750>
 "00000000000000000010110111100111", -- 11750 FREE #<CONS 0 11751>
 "00000000000000000010110111101000", -- 11751 FREE #<CONS 0 11752>
 "00000000000000000010110111101001", -- 11752 FREE #<CONS 0 11753>
 "00000000000000000010110111101010", -- 11753 FREE #<CONS 0 11754>
 "00000000000000000010110111101011", -- 11754 FREE #<CONS 0 11755>
 "00000000000000000010110111101100", -- 11755 FREE #<CONS 0 11756>
 "00000000000000000010110111101101", -- 11756 FREE #<CONS 0 11757>
 "00000000000000000010110111101110", -- 11757 FREE #<CONS 0 11758>
 "00000000000000000010110111101111", -- 11758 FREE #<CONS 0 11759>
 "00000000000000000010110111110000", -- 11759 FREE #<CONS 0 11760>
 "00000000000000000010110111110001", -- 11760 FREE #<CONS 0 11761>
 "00000000000000000010110111110010", -- 11761 FREE #<CONS 0 11762>
 "00000000000000000010110111110011", -- 11762 FREE #<CONS 0 11763>
 "00000000000000000010110111110100", -- 11763 FREE #<CONS 0 11764>
 "00000000000000000010110111110101", -- 11764 FREE #<CONS 0 11765>
 "00000000000000000010110111110110", -- 11765 FREE #<CONS 0 11766>
 "00000000000000000010110111110111", -- 11766 FREE #<CONS 0 11767>
 "00000000000000000010110111111000", -- 11767 FREE #<CONS 0 11768>
 "00000000000000000010110111111001", -- 11768 FREE #<CONS 0 11769>
 "00000000000000000010110111111010", -- 11769 FREE #<CONS 0 11770>
 "00000000000000000010110111111011", -- 11770 FREE #<CONS 0 11771>
 "00000000000000000010110111111100", -- 11771 FREE #<CONS 0 11772>
 "00000000000000000010110111111101", -- 11772 FREE #<CONS 0 11773>
 "00000000000000000010110111111110", -- 11773 FREE #<CONS 0 11774>
 "00000000000000000010110111111111", -- 11774 FREE #<CONS 0 11775>
 "00000000000000000010111000000000", -- 11775 FREE #<CONS 0 11776>
 "00000000000000000010111000000001", -- 11776 FREE #<CONS 0 11777>
 "00000000000000000010111000000010", -- 11777 FREE #<CONS 0 11778>
 "00000000000000000010111000000011", -- 11778 FREE #<CONS 0 11779>
 "00000000000000000010111000000100", -- 11779 FREE #<CONS 0 11780>
 "00000000000000000010111000000101", -- 11780 FREE #<CONS 0 11781>
 "00000000000000000010111000000110", -- 11781 FREE #<CONS 0 11782>
 "00000000000000000010111000000111", -- 11782 FREE #<CONS 0 11783>
 "00000000000000000010111000001000", -- 11783 FREE #<CONS 0 11784>
 "00000000000000000010111000001001", -- 11784 FREE #<CONS 0 11785>
 "00000000000000000010111000001010", -- 11785 FREE #<CONS 0 11786>
 "00000000000000000010111000001011", -- 11786 FREE #<CONS 0 11787>
 "00000000000000000010111000001100", -- 11787 FREE #<CONS 0 11788>
 "00000000000000000010111000001101", -- 11788 FREE #<CONS 0 11789>
 "00000000000000000010111000001110", -- 11789 FREE #<CONS 0 11790>
 "00000000000000000010111000001111", -- 11790 FREE #<CONS 0 11791>
 "00000000000000000010111000010000", -- 11791 FREE #<CONS 0 11792>
 "00000000000000000010111000010001", -- 11792 FREE #<CONS 0 11793>
 "00000000000000000010111000010010", -- 11793 FREE #<CONS 0 11794>
 "00000000000000000010111000010011", -- 11794 FREE #<CONS 0 11795>
 "00000000000000000010111000010100", -- 11795 FREE #<CONS 0 11796>
 "00000000000000000010111000010101", -- 11796 FREE #<CONS 0 11797>
 "00000000000000000010111000010110", -- 11797 FREE #<CONS 0 11798>
 "00000000000000000010111000010111", -- 11798 FREE #<CONS 0 11799>
 "00000000000000000010111000011000", -- 11799 FREE #<CONS 0 11800>
 "00000000000000000010111000011001", -- 11800 FREE #<CONS 0 11801>
 "00000000000000000010111000011010", -- 11801 FREE #<CONS 0 11802>
 "00000000000000000010111000011011", -- 11802 FREE #<CONS 0 11803>
 "00000000000000000010111000011100", -- 11803 FREE #<CONS 0 11804>
 "00000000000000000010111000011101", -- 11804 FREE #<CONS 0 11805>
 "00000000000000000010111000011110", -- 11805 FREE #<CONS 0 11806>
 "00000000000000000010111000011111", -- 11806 FREE #<CONS 0 11807>
 "00000000000000000010111000100000", -- 11807 FREE #<CONS 0 11808>
 "00000000000000000010111000100001", -- 11808 FREE #<CONS 0 11809>
 "00000000000000000010111000100010", -- 11809 FREE #<CONS 0 11810>
 "00000000000000000010111000100011", -- 11810 FREE #<CONS 0 11811>
 "00000000000000000010111000100100", -- 11811 FREE #<CONS 0 11812>
 "00000000000000000010111000100101", -- 11812 FREE #<CONS 0 11813>
 "00000000000000000010111000100110", -- 11813 FREE #<CONS 0 11814>
 "00000000000000000010111000100111", -- 11814 FREE #<CONS 0 11815>
 "00000000000000000010111000101000", -- 11815 FREE #<CONS 0 11816>
 "00000000000000000010111000101001", -- 11816 FREE #<CONS 0 11817>
 "00000000000000000010111000101010", -- 11817 FREE #<CONS 0 11818>
 "00000000000000000010111000101011", -- 11818 FREE #<CONS 0 11819>
 "00000000000000000010111000101100", -- 11819 FREE #<CONS 0 11820>
 "00000000000000000010111000101101", -- 11820 FREE #<CONS 0 11821>
 "00000000000000000010111000101110", -- 11821 FREE #<CONS 0 11822>
 "00000000000000000010111000101111", -- 11822 FREE #<CONS 0 11823>
 "00000000000000000010111000110000", -- 11823 FREE #<CONS 0 11824>
 "00000000000000000010111000110001", -- 11824 FREE #<CONS 0 11825>
 "00000000000000000010111000110010", -- 11825 FREE #<CONS 0 11826>
 "00000000000000000010111000110011", -- 11826 FREE #<CONS 0 11827>
 "00000000000000000010111000110100", -- 11827 FREE #<CONS 0 11828>
 "00000000000000000010111000110101", -- 11828 FREE #<CONS 0 11829>
 "00000000000000000010111000110110", -- 11829 FREE #<CONS 0 11830>
 "00000000000000000010111000110111", -- 11830 FREE #<CONS 0 11831>
 "00000000000000000010111000111000", -- 11831 FREE #<CONS 0 11832>
 "00000000000000000010111000111001", -- 11832 FREE #<CONS 0 11833>
 "00000000000000000010111000111010", -- 11833 FREE #<CONS 0 11834>
 "00000000000000000010111000111011", -- 11834 FREE #<CONS 0 11835>
 "00000000000000000010111000111100", -- 11835 FREE #<CONS 0 11836>
 "00000000000000000010111000111101", -- 11836 FREE #<CONS 0 11837>
 "00000000000000000010111000111110", -- 11837 FREE #<CONS 0 11838>
 "00000000000000000010111000111111", -- 11838 FREE #<CONS 0 11839>
 "00000000000000000010111001000000", -- 11839 FREE #<CONS 0 11840>
 "00000000000000000010111001000001", -- 11840 FREE #<CONS 0 11841>
 "00000000000000000010111001000010", -- 11841 FREE #<CONS 0 11842>
 "00000000000000000010111001000011", -- 11842 FREE #<CONS 0 11843>
 "00000000000000000010111001000100", -- 11843 FREE #<CONS 0 11844>
 "00000000000000000010111001000101", -- 11844 FREE #<CONS 0 11845>
 "00000000000000000010111001000110", -- 11845 FREE #<CONS 0 11846>
 "00000000000000000010111001000111", -- 11846 FREE #<CONS 0 11847>
 "00000000000000000010111001001000", -- 11847 FREE #<CONS 0 11848>
 "00000000000000000010111001001001", -- 11848 FREE #<CONS 0 11849>
 "00000000000000000010111001001010", -- 11849 FREE #<CONS 0 11850>
 "00000000000000000010111001001011", -- 11850 FREE #<CONS 0 11851>
 "00000000000000000010111001001100", -- 11851 FREE #<CONS 0 11852>
 "00000000000000000010111001001101", -- 11852 FREE #<CONS 0 11853>
 "00000000000000000010111001001110", -- 11853 FREE #<CONS 0 11854>
 "00000000000000000010111001001111", -- 11854 FREE #<CONS 0 11855>
 "00000000000000000010111001010000", -- 11855 FREE #<CONS 0 11856>
 "00000000000000000010111001010001", -- 11856 FREE #<CONS 0 11857>
 "00000000000000000010111001010010", -- 11857 FREE #<CONS 0 11858>
 "00000000000000000010111001010011", -- 11858 FREE #<CONS 0 11859>
 "00000000000000000010111001010100", -- 11859 FREE #<CONS 0 11860>
 "00000000000000000010111001010101", -- 11860 FREE #<CONS 0 11861>
 "00000000000000000010111001010110", -- 11861 FREE #<CONS 0 11862>
 "00000000000000000010111001010111", -- 11862 FREE #<CONS 0 11863>
 "00000000000000000010111001011000", -- 11863 FREE #<CONS 0 11864>
 "00000000000000000010111001011001", -- 11864 FREE #<CONS 0 11865>
 "00000000000000000010111001011010", -- 11865 FREE #<CONS 0 11866>
 "00000000000000000010111001011011", -- 11866 FREE #<CONS 0 11867>
 "00000000000000000010111001011100", -- 11867 FREE #<CONS 0 11868>
 "00000000000000000010111001011101", -- 11868 FREE #<CONS 0 11869>
 "00000000000000000010111001011110", -- 11869 FREE #<CONS 0 11870>
 "00000000000000000010111001011111", -- 11870 FREE #<CONS 0 11871>
 "00000000000000000010111001100000", -- 11871 FREE #<CONS 0 11872>
 "00000000000000000010111001100001", -- 11872 FREE #<CONS 0 11873>
 "00000000000000000010111001100010", -- 11873 FREE #<CONS 0 11874>
 "00000000000000000010111001100011", -- 11874 FREE #<CONS 0 11875>
 "00000000000000000010111001100100", -- 11875 FREE #<CONS 0 11876>
 "00000000000000000010111001100101", -- 11876 FREE #<CONS 0 11877>
 "00000000000000000010111001100110", -- 11877 FREE #<CONS 0 11878>
 "00000000000000000010111001100111", -- 11878 FREE #<CONS 0 11879>
 "00000000000000000010111001101000", -- 11879 FREE #<CONS 0 11880>
 "00000000000000000010111001101001", -- 11880 FREE #<CONS 0 11881>
 "00000000000000000010111001101010", -- 11881 FREE #<CONS 0 11882>
 "00000000000000000010111001101011", -- 11882 FREE #<CONS 0 11883>
 "00000000000000000010111001101100", -- 11883 FREE #<CONS 0 11884>
 "00000000000000000010111001101101", -- 11884 FREE #<CONS 0 11885>
 "00000000000000000010111001101110", -- 11885 FREE #<CONS 0 11886>
 "00000000000000000010111001101111", -- 11886 FREE #<CONS 0 11887>
 "00000000000000000010111001110000", -- 11887 FREE #<CONS 0 11888>
 "00000000000000000010111001110001", -- 11888 FREE #<CONS 0 11889>
 "00000000000000000010111001110010", -- 11889 FREE #<CONS 0 11890>
 "00000000000000000010111001110011", -- 11890 FREE #<CONS 0 11891>
 "00000000000000000010111001110100", -- 11891 FREE #<CONS 0 11892>
 "00000000000000000010111001110101", -- 11892 FREE #<CONS 0 11893>
 "00000000000000000010111001110110", -- 11893 FREE #<CONS 0 11894>
 "00000000000000000010111001110111", -- 11894 FREE #<CONS 0 11895>
 "00000000000000000010111001111000", -- 11895 FREE #<CONS 0 11896>
 "00000000000000000010111001111001", -- 11896 FREE #<CONS 0 11897>
 "00000000000000000010111001111010", -- 11897 FREE #<CONS 0 11898>
 "00000000000000000010111001111011", -- 11898 FREE #<CONS 0 11899>
 "00000000000000000010111001111100", -- 11899 FREE #<CONS 0 11900>
 "00000000000000000010111001111101", -- 11900 FREE #<CONS 0 11901>
 "00000000000000000010111001111110", -- 11901 FREE #<CONS 0 11902>
 "00000000000000000010111001111111", -- 11902 FREE #<CONS 0 11903>
 "00000000000000000010111010000000", -- 11903 FREE #<CONS 0 11904>
 "00000000000000000010111010000001", -- 11904 FREE #<CONS 0 11905>
 "00000000000000000010111010000010", -- 11905 FREE #<CONS 0 11906>
 "00000000000000000010111010000011", -- 11906 FREE #<CONS 0 11907>
 "00000000000000000010111010000100", -- 11907 FREE #<CONS 0 11908>
 "00000000000000000010111010000101", -- 11908 FREE #<CONS 0 11909>
 "00000000000000000010111010000110", -- 11909 FREE #<CONS 0 11910>
 "00000000000000000010111010000111", -- 11910 FREE #<CONS 0 11911>
 "00000000000000000010111010001000", -- 11911 FREE #<CONS 0 11912>
 "00000000000000000010111010001001", -- 11912 FREE #<CONS 0 11913>
 "00000000000000000010111010001010", -- 11913 FREE #<CONS 0 11914>
 "00000000000000000010111010001011", -- 11914 FREE #<CONS 0 11915>
 "00000000000000000010111010001100", -- 11915 FREE #<CONS 0 11916>
 "00000000000000000010111010001101", -- 11916 FREE #<CONS 0 11917>
 "00000000000000000010111010001110", -- 11917 FREE #<CONS 0 11918>
 "00000000000000000010111010001111", -- 11918 FREE #<CONS 0 11919>
 "00000000000000000010111010010000", -- 11919 FREE #<CONS 0 11920>
 "00000000000000000010111010010001", -- 11920 FREE #<CONS 0 11921>
 "00000000000000000010111010010010", -- 11921 FREE #<CONS 0 11922>
 "00000000000000000010111010010011", -- 11922 FREE #<CONS 0 11923>
 "00000000000000000010111010010100", -- 11923 FREE #<CONS 0 11924>
 "00000000000000000010111010010101", -- 11924 FREE #<CONS 0 11925>
 "00000000000000000010111010010110", -- 11925 FREE #<CONS 0 11926>
 "00000000000000000010111010010111", -- 11926 FREE #<CONS 0 11927>
 "00000000000000000010111010011000", -- 11927 FREE #<CONS 0 11928>
 "00000000000000000010111010011001", -- 11928 FREE #<CONS 0 11929>
 "00000000000000000010111010011010", -- 11929 FREE #<CONS 0 11930>
 "00000000000000000010111010011011", -- 11930 FREE #<CONS 0 11931>
 "00000000000000000010111010011100", -- 11931 FREE #<CONS 0 11932>
 "00000000000000000010111010011101", -- 11932 FREE #<CONS 0 11933>
 "00000000000000000010111010011110", -- 11933 FREE #<CONS 0 11934>
 "00000000000000000010111010011111", -- 11934 FREE #<CONS 0 11935>
 "00000000000000000010111010100000", -- 11935 FREE #<CONS 0 11936>
 "00000000000000000010111010100001", -- 11936 FREE #<CONS 0 11937>
 "00000000000000000010111010100010", -- 11937 FREE #<CONS 0 11938>
 "00000000000000000010111010100011", -- 11938 FREE #<CONS 0 11939>
 "00000000000000000010111010100100", -- 11939 FREE #<CONS 0 11940>
 "00000000000000000010111010100101", -- 11940 FREE #<CONS 0 11941>
 "00000000000000000010111010100110", -- 11941 FREE #<CONS 0 11942>
 "00000000000000000010111010100111", -- 11942 FREE #<CONS 0 11943>
 "00000000000000000010111010101000", -- 11943 FREE #<CONS 0 11944>
 "00000000000000000010111010101001", -- 11944 FREE #<CONS 0 11945>
 "00000000000000000010111010101010", -- 11945 FREE #<CONS 0 11946>
 "00000000000000000010111010101011", -- 11946 FREE #<CONS 0 11947>
 "00000000000000000010111010101100", -- 11947 FREE #<CONS 0 11948>
 "00000000000000000010111010101101", -- 11948 FREE #<CONS 0 11949>
 "00000000000000000010111010101110", -- 11949 FREE #<CONS 0 11950>
 "00000000000000000010111010101111", -- 11950 FREE #<CONS 0 11951>
 "00000000000000000010111010110000", -- 11951 FREE #<CONS 0 11952>
 "00000000000000000010111010110001", -- 11952 FREE #<CONS 0 11953>
 "00000000000000000010111010110010", -- 11953 FREE #<CONS 0 11954>
 "00000000000000000010111010110011", -- 11954 FREE #<CONS 0 11955>
 "00000000000000000010111010110100", -- 11955 FREE #<CONS 0 11956>
 "00000000000000000010111010110101", -- 11956 FREE #<CONS 0 11957>
 "00000000000000000010111010110110", -- 11957 FREE #<CONS 0 11958>
 "00000000000000000010111010110111", -- 11958 FREE #<CONS 0 11959>
 "00000000000000000010111010111000", -- 11959 FREE #<CONS 0 11960>
 "00000000000000000010111010111001", -- 11960 FREE #<CONS 0 11961>
 "00000000000000000010111010111010", -- 11961 FREE #<CONS 0 11962>
 "00000000000000000010111010111011", -- 11962 FREE #<CONS 0 11963>
 "00000000000000000010111010111100", -- 11963 FREE #<CONS 0 11964>
 "00000000000000000010111010111101", -- 11964 FREE #<CONS 0 11965>
 "00000000000000000010111010111110", -- 11965 FREE #<CONS 0 11966>
 "00000000000000000010111010111111", -- 11966 FREE #<CONS 0 11967>
 "00000000000000000010111011000000", -- 11967 FREE #<CONS 0 11968>
 "00000000000000000010111011000001", -- 11968 FREE #<CONS 0 11969>
 "00000000000000000010111011000010", -- 11969 FREE #<CONS 0 11970>
 "00000000000000000010111011000011", -- 11970 FREE #<CONS 0 11971>
 "00000000000000000010111011000100", -- 11971 FREE #<CONS 0 11972>
 "00000000000000000010111011000101", -- 11972 FREE #<CONS 0 11973>
 "00000000000000000010111011000110", -- 11973 FREE #<CONS 0 11974>
 "00000000000000000010111011000111", -- 11974 FREE #<CONS 0 11975>
 "00000000000000000010111011001000", -- 11975 FREE #<CONS 0 11976>
 "00000000000000000010111011001001", -- 11976 FREE #<CONS 0 11977>
 "00000000000000000010111011001010", -- 11977 FREE #<CONS 0 11978>
 "00000000000000000010111011001011", -- 11978 FREE #<CONS 0 11979>
 "00000000000000000010111011001100", -- 11979 FREE #<CONS 0 11980>
 "00000000000000000010111011001101", -- 11980 FREE #<CONS 0 11981>
 "00000000000000000010111011001110", -- 11981 FREE #<CONS 0 11982>
 "00000000000000000010111011001111", -- 11982 FREE #<CONS 0 11983>
 "00000000000000000010111011010000", -- 11983 FREE #<CONS 0 11984>
 "00000000000000000010111011010001", -- 11984 FREE #<CONS 0 11985>
 "00000000000000000010111011010010", -- 11985 FREE #<CONS 0 11986>
 "00000000000000000010111011010011", -- 11986 FREE #<CONS 0 11987>
 "00000000000000000010111011010100", -- 11987 FREE #<CONS 0 11988>
 "00000000000000000010111011010101", -- 11988 FREE #<CONS 0 11989>
 "00000000000000000010111011010110", -- 11989 FREE #<CONS 0 11990>
 "00000000000000000010111011010111", -- 11990 FREE #<CONS 0 11991>
 "00000000000000000010111011011000", -- 11991 FREE #<CONS 0 11992>
 "00000000000000000010111011011001", -- 11992 FREE #<CONS 0 11993>
 "00000000000000000010111011011010", -- 11993 FREE #<CONS 0 11994>
 "00000000000000000010111011011011", -- 11994 FREE #<CONS 0 11995>
 "00000000000000000010111011011100", -- 11995 FREE #<CONS 0 11996>
 "00000000000000000010111011011101", -- 11996 FREE #<CONS 0 11997>
 "00000000000000000010111011011110", -- 11997 FREE #<CONS 0 11998>
 "00000000000000000010111011011111", -- 11998 FREE #<CONS 0 11999>
 "00000000000000000010111011100000", -- 11999 FREE #<CONS 0 12000>
 "00000000000000000010111011100001", -- 12000 FREE #<CONS 0 12001>
 "00000000000000000010111011100010", -- 12001 FREE #<CONS 0 12002>
 "00000000000000000010111011100011", -- 12002 FREE #<CONS 0 12003>
 "00000000000000000010111011100100", -- 12003 FREE #<CONS 0 12004>
 "00000000000000000010111011100101", -- 12004 FREE #<CONS 0 12005>
 "00000000000000000010111011100110", -- 12005 FREE #<CONS 0 12006>
 "00000000000000000010111011100111", -- 12006 FREE #<CONS 0 12007>
 "00000000000000000010111011101000", -- 12007 FREE #<CONS 0 12008>
 "00000000000000000010111011101001", -- 12008 FREE #<CONS 0 12009>
 "00000000000000000010111011101010", -- 12009 FREE #<CONS 0 12010>
 "00000000000000000010111011101011", -- 12010 FREE #<CONS 0 12011>
 "00000000000000000010111011101100", -- 12011 FREE #<CONS 0 12012>
 "00000000000000000010111011101101", -- 12012 FREE #<CONS 0 12013>
 "00000000000000000010111011101110", -- 12013 FREE #<CONS 0 12014>
 "00000000000000000010111011101111", -- 12014 FREE #<CONS 0 12015>
 "00000000000000000010111011110000", -- 12015 FREE #<CONS 0 12016>
 "00000000000000000010111011110001", -- 12016 FREE #<CONS 0 12017>
 "00000000000000000010111011110010", -- 12017 FREE #<CONS 0 12018>
 "00000000000000000010111011110011", -- 12018 FREE #<CONS 0 12019>
 "00000000000000000010111011110100", -- 12019 FREE #<CONS 0 12020>
 "00000000000000000010111011110101", -- 12020 FREE #<CONS 0 12021>
 "00000000000000000010111011110110", -- 12021 FREE #<CONS 0 12022>
 "00000000000000000010111011110111", -- 12022 FREE #<CONS 0 12023>
 "00000000000000000010111011111000", -- 12023 FREE #<CONS 0 12024>
 "00000000000000000010111011111001", -- 12024 FREE #<CONS 0 12025>
 "00000000000000000010111011111010", -- 12025 FREE #<CONS 0 12026>
 "00000000000000000010111011111011", -- 12026 FREE #<CONS 0 12027>
 "00000000000000000010111011111100", -- 12027 FREE #<CONS 0 12028>
 "00000000000000000010111011111101", -- 12028 FREE #<CONS 0 12029>
 "00000000000000000010111011111110", -- 12029 FREE #<CONS 0 12030>
 "00000000000000000010111011111111", -- 12030 FREE #<CONS 0 12031>
 "00000000000000000010111100000000", -- 12031 FREE #<CONS 0 12032>
 "00000000000000000010111100000001", -- 12032 FREE #<CONS 0 12033>
 "00000000000000000010111100000010", -- 12033 FREE #<CONS 0 12034>
 "00000000000000000010111100000011", -- 12034 FREE #<CONS 0 12035>
 "00000000000000000010111100000100", -- 12035 FREE #<CONS 0 12036>
 "00000000000000000010111100000101", -- 12036 FREE #<CONS 0 12037>
 "00000000000000000010111100000110", -- 12037 FREE #<CONS 0 12038>
 "00000000000000000010111100000111", -- 12038 FREE #<CONS 0 12039>
 "00000000000000000010111100001000", -- 12039 FREE #<CONS 0 12040>
 "00000000000000000010111100001001", -- 12040 FREE #<CONS 0 12041>
 "00000000000000000010111100001010", -- 12041 FREE #<CONS 0 12042>
 "00000000000000000010111100001011", -- 12042 FREE #<CONS 0 12043>
 "00000000000000000010111100001100", -- 12043 FREE #<CONS 0 12044>
 "00000000000000000010111100001101", -- 12044 FREE #<CONS 0 12045>
 "00000000000000000010111100001110", -- 12045 FREE #<CONS 0 12046>
 "00000000000000000010111100001111", -- 12046 FREE #<CONS 0 12047>
 "00000000000000000010111100010000", -- 12047 FREE #<CONS 0 12048>
 "00000000000000000010111100010001", -- 12048 FREE #<CONS 0 12049>
 "00000000000000000010111100010010", -- 12049 FREE #<CONS 0 12050>
 "00000000000000000010111100010011", -- 12050 FREE #<CONS 0 12051>
 "00000000000000000010111100010100", -- 12051 FREE #<CONS 0 12052>
 "00000000000000000010111100010101", -- 12052 FREE #<CONS 0 12053>
 "00000000000000000010111100010110", -- 12053 FREE #<CONS 0 12054>
 "00000000000000000010111100010111", -- 12054 FREE #<CONS 0 12055>
 "00000000000000000010111100011000", -- 12055 FREE #<CONS 0 12056>
 "00000000000000000010111100011001", -- 12056 FREE #<CONS 0 12057>
 "00000000000000000010111100011010", -- 12057 FREE #<CONS 0 12058>
 "00000000000000000010111100011011", -- 12058 FREE #<CONS 0 12059>
 "00000000000000000010111100011100", -- 12059 FREE #<CONS 0 12060>
 "00000000000000000010111100011101", -- 12060 FREE #<CONS 0 12061>
 "00000000000000000010111100011110", -- 12061 FREE #<CONS 0 12062>
 "00000000000000000010111100011111", -- 12062 FREE #<CONS 0 12063>
 "00000000000000000010111100100000", -- 12063 FREE #<CONS 0 12064>
 "00000000000000000010111100100001", -- 12064 FREE #<CONS 0 12065>
 "00000000000000000010111100100010", -- 12065 FREE #<CONS 0 12066>
 "00000000000000000010111100100011", -- 12066 FREE #<CONS 0 12067>
 "00000000000000000010111100100100", -- 12067 FREE #<CONS 0 12068>
 "00000000000000000010111100100101", -- 12068 FREE #<CONS 0 12069>
 "00000000000000000010111100100110", -- 12069 FREE #<CONS 0 12070>
 "00000000000000000010111100100111", -- 12070 FREE #<CONS 0 12071>
 "00000000000000000010111100101000", -- 12071 FREE #<CONS 0 12072>
 "00000000000000000010111100101001", -- 12072 FREE #<CONS 0 12073>
 "00000000000000000010111100101010", -- 12073 FREE #<CONS 0 12074>
 "00000000000000000010111100101011", -- 12074 FREE #<CONS 0 12075>
 "00000000000000000010111100101100", -- 12075 FREE #<CONS 0 12076>
 "00000000000000000010111100101101", -- 12076 FREE #<CONS 0 12077>
 "00000000000000000010111100101110", -- 12077 FREE #<CONS 0 12078>
 "00000000000000000010111100101111", -- 12078 FREE #<CONS 0 12079>
 "00000000000000000010111100110000", -- 12079 FREE #<CONS 0 12080>
 "00000000000000000010111100110001", -- 12080 FREE #<CONS 0 12081>
 "00000000000000000010111100110010", -- 12081 FREE #<CONS 0 12082>
 "00000000000000000010111100110011", -- 12082 FREE #<CONS 0 12083>
 "00000000000000000010111100110100", -- 12083 FREE #<CONS 0 12084>
 "00000000000000000010111100110101", -- 12084 FREE #<CONS 0 12085>
 "00000000000000000010111100110110", -- 12085 FREE #<CONS 0 12086>
 "00000000000000000010111100110111", -- 12086 FREE #<CONS 0 12087>
 "00000000000000000010111100111000", -- 12087 FREE #<CONS 0 12088>
 "00000000000000000010111100111001", -- 12088 FREE #<CONS 0 12089>
 "00000000000000000010111100111010", -- 12089 FREE #<CONS 0 12090>
 "00000000000000000010111100111011", -- 12090 FREE #<CONS 0 12091>
 "00000000000000000010111100111100", -- 12091 FREE #<CONS 0 12092>
 "00000000000000000010111100111101", -- 12092 FREE #<CONS 0 12093>
 "00000000000000000010111100111110", -- 12093 FREE #<CONS 0 12094>
 "00000000000000000010111100111111", -- 12094 FREE #<CONS 0 12095>
 "00000000000000000010111101000000", -- 12095 FREE #<CONS 0 12096>
 "00000000000000000010111101000001", -- 12096 FREE #<CONS 0 12097>
 "00000000000000000010111101000010", -- 12097 FREE #<CONS 0 12098>
 "00000000000000000010111101000011", -- 12098 FREE #<CONS 0 12099>
 "00000000000000000010111101000100", -- 12099 FREE #<CONS 0 12100>
 "00000000000000000010111101000101", -- 12100 FREE #<CONS 0 12101>
 "00000000000000000010111101000110", -- 12101 FREE #<CONS 0 12102>
 "00000000000000000010111101000111", -- 12102 FREE #<CONS 0 12103>
 "00000000000000000010111101001000", -- 12103 FREE #<CONS 0 12104>
 "00000000000000000010111101001001", -- 12104 FREE #<CONS 0 12105>
 "00000000000000000010111101001010", -- 12105 FREE #<CONS 0 12106>
 "00000000000000000010111101001011", -- 12106 FREE #<CONS 0 12107>
 "00000000000000000010111101001100", -- 12107 FREE #<CONS 0 12108>
 "00000000000000000010111101001101", -- 12108 FREE #<CONS 0 12109>
 "00000000000000000010111101001110", -- 12109 FREE #<CONS 0 12110>
 "00000000000000000010111101001111", -- 12110 FREE #<CONS 0 12111>
 "00000000000000000010111101010000", -- 12111 FREE #<CONS 0 12112>
 "00000000000000000010111101010001", -- 12112 FREE #<CONS 0 12113>
 "00000000000000000010111101010010", -- 12113 FREE #<CONS 0 12114>
 "00000000000000000010111101010011", -- 12114 FREE #<CONS 0 12115>
 "00000000000000000010111101010100", -- 12115 FREE #<CONS 0 12116>
 "00000000000000000010111101010101", -- 12116 FREE #<CONS 0 12117>
 "00000000000000000010111101010110", -- 12117 FREE #<CONS 0 12118>
 "00000000000000000010111101010111", -- 12118 FREE #<CONS 0 12119>
 "00000000000000000010111101011000", -- 12119 FREE #<CONS 0 12120>
 "00000000000000000010111101011001", -- 12120 FREE #<CONS 0 12121>
 "00000000000000000010111101011010", -- 12121 FREE #<CONS 0 12122>
 "00000000000000000010111101011011", -- 12122 FREE #<CONS 0 12123>
 "00000000000000000010111101011100", -- 12123 FREE #<CONS 0 12124>
 "00000000000000000010111101011101", -- 12124 FREE #<CONS 0 12125>
 "00000000000000000010111101011110", -- 12125 FREE #<CONS 0 12126>
 "00000000000000000010111101011111", -- 12126 FREE #<CONS 0 12127>
 "00000000000000000010111101100000", -- 12127 FREE #<CONS 0 12128>
 "00000000000000000010111101100001", -- 12128 FREE #<CONS 0 12129>
 "00000000000000000010111101100010", -- 12129 FREE #<CONS 0 12130>
 "00000000000000000010111101100011", -- 12130 FREE #<CONS 0 12131>
 "00000000000000000010111101100100", -- 12131 FREE #<CONS 0 12132>
 "00000000000000000010111101100101", -- 12132 FREE #<CONS 0 12133>
 "00000000000000000010111101100110", -- 12133 FREE #<CONS 0 12134>
 "00000000000000000010111101100111", -- 12134 FREE #<CONS 0 12135>
 "00000000000000000010111101101000", -- 12135 FREE #<CONS 0 12136>
 "00000000000000000010111101101001", -- 12136 FREE #<CONS 0 12137>
 "00000000000000000010111101101010", -- 12137 FREE #<CONS 0 12138>
 "00000000000000000010111101101011", -- 12138 FREE #<CONS 0 12139>
 "00000000000000000010111101101100", -- 12139 FREE #<CONS 0 12140>
 "00000000000000000010111101101101", -- 12140 FREE #<CONS 0 12141>
 "00000000000000000010111101101110", -- 12141 FREE #<CONS 0 12142>
 "00000000000000000010111101101111", -- 12142 FREE #<CONS 0 12143>
 "00000000000000000010111101110000", -- 12143 FREE #<CONS 0 12144>
 "00000000000000000010111101110001", -- 12144 FREE #<CONS 0 12145>
 "00000000000000000010111101110010", -- 12145 FREE #<CONS 0 12146>
 "00000000000000000010111101110011", -- 12146 FREE #<CONS 0 12147>
 "00000000000000000010111101110100", -- 12147 FREE #<CONS 0 12148>
 "00000000000000000010111101110101", -- 12148 FREE #<CONS 0 12149>
 "00000000000000000010111101110110", -- 12149 FREE #<CONS 0 12150>
 "00000000000000000010111101110111", -- 12150 FREE #<CONS 0 12151>
 "00000000000000000010111101111000", -- 12151 FREE #<CONS 0 12152>
 "00000000000000000010111101111001", -- 12152 FREE #<CONS 0 12153>
 "00000000000000000010111101111010", -- 12153 FREE #<CONS 0 12154>
 "00000000000000000010111101111011", -- 12154 FREE #<CONS 0 12155>
 "00000000000000000010111101111100", -- 12155 FREE #<CONS 0 12156>
 "00000000000000000010111101111101", -- 12156 FREE #<CONS 0 12157>
 "00000000000000000010111101111110", -- 12157 FREE #<CONS 0 12158>
 "00000000000000000010111101111111", -- 12158 FREE #<CONS 0 12159>
 "00000000000000000010111110000000", -- 12159 FREE #<CONS 0 12160>
 "00000000000000000010111110000001", -- 12160 FREE #<CONS 0 12161>
 "00000000000000000010111110000010", -- 12161 FREE #<CONS 0 12162>
 "00000000000000000010111110000011", -- 12162 FREE #<CONS 0 12163>
 "00000000000000000010111110000100", -- 12163 FREE #<CONS 0 12164>
 "00000000000000000010111110000101", -- 12164 FREE #<CONS 0 12165>
 "00000000000000000010111110000110", -- 12165 FREE #<CONS 0 12166>
 "00000000000000000010111110000111", -- 12166 FREE #<CONS 0 12167>
 "00000000000000000010111110001000", -- 12167 FREE #<CONS 0 12168>
 "00000000000000000010111110001001", -- 12168 FREE #<CONS 0 12169>
 "00000000000000000010111110001010", -- 12169 FREE #<CONS 0 12170>
 "00000000000000000010111110001011", -- 12170 FREE #<CONS 0 12171>
 "00000000000000000010111110001100", -- 12171 FREE #<CONS 0 12172>
 "00000000000000000010111110001101", -- 12172 FREE #<CONS 0 12173>
 "00000000000000000010111110001110", -- 12173 FREE #<CONS 0 12174>
 "00000000000000000010111110001111", -- 12174 FREE #<CONS 0 12175>
 "00000000000000000010111110010000", -- 12175 FREE #<CONS 0 12176>
 "00000000000000000010111110010001", -- 12176 FREE #<CONS 0 12177>
 "00000000000000000010111110010010", -- 12177 FREE #<CONS 0 12178>
 "00000000000000000010111110010011", -- 12178 FREE #<CONS 0 12179>
 "00000000000000000010111110010100", -- 12179 FREE #<CONS 0 12180>
 "00000000000000000010111110010101", -- 12180 FREE #<CONS 0 12181>
 "00000000000000000010111110010110", -- 12181 FREE #<CONS 0 12182>
 "00000000000000000010111110010111", -- 12182 FREE #<CONS 0 12183>
 "00000000000000000010111110011000", -- 12183 FREE #<CONS 0 12184>
 "00000000000000000010111110011001", -- 12184 FREE #<CONS 0 12185>
 "00000000000000000010111110011010", -- 12185 FREE #<CONS 0 12186>
 "00000000000000000010111110011011", -- 12186 FREE #<CONS 0 12187>
 "00000000000000000010111110011100", -- 12187 FREE #<CONS 0 12188>
 "00000000000000000010111110011101", -- 12188 FREE #<CONS 0 12189>
 "00000000000000000010111110011110", -- 12189 FREE #<CONS 0 12190>
 "00000000000000000010111110011111", -- 12190 FREE #<CONS 0 12191>
 "00000000000000000010111110100000", -- 12191 FREE #<CONS 0 12192>
 "00000000000000000010111110100001", -- 12192 FREE #<CONS 0 12193>
 "00000000000000000010111110100010", -- 12193 FREE #<CONS 0 12194>
 "00000000000000000010111110100011", -- 12194 FREE #<CONS 0 12195>
 "00000000000000000010111110100100", -- 12195 FREE #<CONS 0 12196>
 "00000000000000000010111110100101", -- 12196 FREE #<CONS 0 12197>
 "00000000000000000010111110100110", -- 12197 FREE #<CONS 0 12198>
 "00000000000000000010111110100111", -- 12198 FREE #<CONS 0 12199>
 "00000000000000000010111110101000", -- 12199 FREE #<CONS 0 12200>
 "00000000000000000010111110101001", -- 12200 FREE #<CONS 0 12201>
 "00000000000000000010111110101010", -- 12201 FREE #<CONS 0 12202>
 "00000000000000000010111110101011", -- 12202 FREE #<CONS 0 12203>
 "00000000000000000010111110101100", -- 12203 FREE #<CONS 0 12204>
 "00000000000000000010111110101101", -- 12204 FREE #<CONS 0 12205>
 "00000000000000000010111110101110", -- 12205 FREE #<CONS 0 12206>
 "00000000000000000010111110101111", -- 12206 FREE #<CONS 0 12207>
 "00000000000000000010111110110000", -- 12207 FREE #<CONS 0 12208>
 "00000000000000000010111110110001", -- 12208 FREE #<CONS 0 12209>
 "00000000000000000010111110110010", -- 12209 FREE #<CONS 0 12210>
 "00000000000000000010111110110011", -- 12210 FREE #<CONS 0 12211>
 "00000000000000000010111110110100", -- 12211 FREE #<CONS 0 12212>
 "00000000000000000010111110110101", -- 12212 FREE #<CONS 0 12213>
 "00000000000000000010111110110110", -- 12213 FREE #<CONS 0 12214>
 "00000000000000000010111110110111", -- 12214 FREE #<CONS 0 12215>
 "00000000000000000010111110111000", -- 12215 FREE #<CONS 0 12216>
 "00000000000000000010111110111001", -- 12216 FREE #<CONS 0 12217>
 "00000000000000000010111110111010", -- 12217 FREE #<CONS 0 12218>
 "00000000000000000010111110111011", -- 12218 FREE #<CONS 0 12219>
 "00000000000000000010111110111100", -- 12219 FREE #<CONS 0 12220>
 "00000000000000000010111110111101", -- 12220 FREE #<CONS 0 12221>
 "00000000000000000010111110111110", -- 12221 FREE #<CONS 0 12222>
 "00000000000000000010111110111111", -- 12222 FREE #<CONS 0 12223>
 "00000000000000000010111111000000", -- 12223 FREE #<CONS 0 12224>
 "00000000000000000010111111000001", -- 12224 FREE #<CONS 0 12225>
 "00000000000000000010111111000010", -- 12225 FREE #<CONS 0 12226>
 "00000000000000000010111111000011", -- 12226 FREE #<CONS 0 12227>
 "00000000000000000010111111000100", -- 12227 FREE #<CONS 0 12228>
 "00000000000000000010111111000101", -- 12228 FREE #<CONS 0 12229>
 "00000000000000000010111111000110", -- 12229 FREE #<CONS 0 12230>
 "00000000000000000010111111000111", -- 12230 FREE #<CONS 0 12231>
 "00000000000000000010111111001000", -- 12231 FREE #<CONS 0 12232>
 "00000000000000000010111111001001", -- 12232 FREE #<CONS 0 12233>
 "00000000000000000010111111001010", -- 12233 FREE #<CONS 0 12234>
 "00000000000000000010111111001011", -- 12234 FREE #<CONS 0 12235>
 "00000000000000000010111111001100", -- 12235 FREE #<CONS 0 12236>
 "00000000000000000010111111001101", -- 12236 FREE #<CONS 0 12237>
 "00000000000000000010111111001110", -- 12237 FREE #<CONS 0 12238>
 "00000000000000000010111111001111", -- 12238 FREE #<CONS 0 12239>
 "00000000000000000010111111010000", -- 12239 FREE #<CONS 0 12240>
 "00000000000000000010111111010001", -- 12240 FREE #<CONS 0 12241>
 "00000000000000000010111111010010", -- 12241 FREE #<CONS 0 12242>
 "00000000000000000010111111010011", -- 12242 FREE #<CONS 0 12243>
 "00000000000000000010111111010100", -- 12243 FREE #<CONS 0 12244>
 "00000000000000000010111111010101", -- 12244 FREE #<CONS 0 12245>
 "00000000000000000010111111010110", -- 12245 FREE #<CONS 0 12246>
 "00000000000000000010111111010111", -- 12246 FREE #<CONS 0 12247>
 "00000000000000000010111111011000", -- 12247 FREE #<CONS 0 12248>
 "00000000000000000010111111011001", -- 12248 FREE #<CONS 0 12249>
 "00000000000000000010111111011010", -- 12249 FREE #<CONS 0 12250>
 "00000000000000000010111111011011", -- 12250 FREE #<CONS 0 12251>
 "00000000000000000010111111011100", -- 12251 FREE #<CONS 0 12252>
 "00000000000000000010111111011101", -- 12252 FREE #<CONS 0 12253>
 "00000000000000000010111111011110", -- 12253 FREE #<CONS 0 12254>
 "00000000000000000010111111011111", -- 12254 FREE #<CONS 0 12255>
 "00000000000000000010111111100000", -- 12255 FREE #<CONS 0 12256>
 "00000000000000000010111111100001", -- 12256 FREE #<CONS 0 12257>
 "00000000000000000010111111100010", -- 12257 FREE #<CONS 0 12258>
 "00000000000000000010111111100011", -- 12258 FREE #<CONS 0 12259>
 "00000000000000000010111111100100", -- 12259 FREE #<CONS 0 12260>
 "00000000000000000010111111100101", -- 12260 FREE #<CONS 0 12261>
 "00000000000000000010111111100110", -- 12261 FREE #<CONS 0 12262>
 "00000000000000000010111111100111", -- 12262 FREE #<CONS 0 12263>
 "00000000000000000010111111101000", -- 12263 FREE #<CONS 0 12264>
 "00000000000000000010111111101001", -- 12264 FREE #<CONS 0 12265>
 "00000000000000000010111111101010", -- 12265 FREE #<CONS 0 12266>
 "00000000000000000010111111101011", -- 12266 FREE #<CONS 0 12267>
 "00000000000000000010111111101100", -- 12267 FREE #<CONS 0 12268>
 "00000000000000000010111111101101", -- 12268 FREE #<CONS 0 12269>
 "00000000000000000010111111101110", -- 12269 FREE #<CONS 0 12270>
 "00000000000000000010111111101111", -- 12270 FREE #<CONS 0 12271>
 "00000000000000000010111111110000", -- 12271 FREE #<CONS 0 12272>
 "00000000000000000010111111110001", -- 12272 FREE #<CONS 0 12273>
 "00000000000000000010111111110010", -- 12273 FREE #<CONS 0 12274>
 "00000000000000000010111111110011", -- 12274 FREE #<CONS 0 12275>
 "00000000000000000010111111110100", -- 12275 FREE #<CONS 0 12276>
 "00000000000000000010111111110101", -- 12276 FREE #<CONS 0 12277>
 "00000000000000000010111111110110", -- 12277 FREE #<CONS 0 12278>
 "00000000000000000010111111110111", -- 12278 FREE #<CONS 0 12279>
 "00000000000000000010111111111000", -- 12279 FREE #<CONS 0 12280>
 "00000000000000000010111111111001", -- 12280 FREE #<CONS 0 12281>
 "00000000000000000010111111111010", -- 12281 FREE #<CONS 0 12282>
 "00000000000000000010111111111011", -- 12282 FREE #<CONS 0 12283>
 "00000000000000000010111111111100", -- 12283 FREE #<CONS 0 12284>
 "00000000000000000010111111111101", -- 12284 FREE #<CONS 0 12285>
 "00000000000000000010111111111110", -- 12285 FREE #<CONS 0 12286>
 "00000000000000000010111111111111", -- 12286 FREE #<CONS 0 12287>
 "00000000000000000011000000000000", -- 12287 FREE #<CONS 0 12288>
 "00000000000000000011000000000001", -- 12288 FREE #<CONS 0 12289>
 "00000000000000000011000000000010", -- 12289 FREE #<CONS 0 12290>
 "00000000000000000011000000000011", -- 12290 FREE #<CONS 0 12291>
 "00000000000000000011000000000100", -- 12291 FREE #<CONS 0 12292>
 "00000000000000000011000000000101", -- 12292 FREE #<CONS 0 12293>
 "00000000000000000011000000000110", -- 12293 FREE #<CONS 0 12294>
 "00000000000000000011000000000111", -- 12294 FREE #<CONS 0 12295>
 "00000000000000000011000000001000", -- 12295 FREE #<CONS 0 12296>
 "00000000000000000011000000001001", -- 12296 FREE #<CONS 0 12297>
 "00000000000000000011000000001010", -- 12297 FREE #<CONS 0 12298>
 "00000000000000000011000000001011", -- 12298 FREE #<CONS 0 12299>
 "00000000000000000011000000001100", -- 12299 FREE #<CONS 0 12300>
 "00000000000000000011000000001101", -- 12300 FREE #<CONS 0 12301>
 "00000000000000000011000000001110", -- 12301 FREE #<CONS 0 12302>
 "00000000000000000011000000001111", -- 12302 FREE #<CONS 0 12303>
 "00000000000000000011000000010000", -- 12303 FREE #<CONS 0 12304>
 "00000000000000000011000000010001", -- 12304 FREE #<CONS 0 12305>
 "00000000000000000011000000010010", -- 12305 FREE #<CONS 0 12306>
 "00000000000000000011000000010011", -- 12306 FREE #<CONS 0 12307>
 "00000000000000000011000000010100", -- 12307 FREE #<CONS 0 12308>
 "00000000000000000011000000010101", -- 12308 FREE #<CONS 0 12309>
 "00000000000000000011000000010110", -- 12309 FREE #<CONS 0 12310>
 "00000000000000000011000000010111", -- 12310 FREE #<CONS 0 12311>
 "00000000000000000011000000011000", -- 12311 FREE #<CONS 0 12312>
 "00000000000000000011000000011001", -- 12312 FREE #<CONS 0 12313>
 "00000000000000000011000000011010", -- 12313 FREE #<CONS 0 12314>
 "00000000000000000011000000011011", -- 12314 FREE #<CONS 0 12315>
 "00000000000000000011000000011100", -- 12315 FREE #<CONS 0 12316>
 "00000000000000000011000000011101", -- 12316 FREE #<CONS 0 12317>
 "00000000000000000011000000011110", -- 12317 FREE #<CONS 0 12318>
 "00000000000000000011000000011111", -- 12318 FREE #<CONS 0 12319>
 "00000000000000000011000000100000", -- 12319 FREE #<CONS 0 12320>
 "00000000000000000011000000100001", -- 12320 FREE #<CONS 0 12321>
 "00000000000000000011000000100010", -- 12321 FREE #<CONS 0 12322>
 "00000000000000000011000000100011", -- 12322 FREE #<CONS 0 12323>
 "00000000000000000011000000100100", -- 12323 FREE #<CONS 0 12324>
 "00000000000000000011000000100101", -- 12324 FREE #<CONS 0 12325>
 "00000000000000000011000000100110", -- 12325 FREE #<CONS 0 12326>
 "00000000000000000011000000100111", -- 12326 FREE #<CONS 0 12327>
 "00000000000000000011000000101000", -- 12327 FREE #<CONS 0 12328>
 "00000000000000000011000000101001", -- 12328 FREE #<CONS 0 12329>
 "00000000000000000011000000101010", -- 12329 FREE #<CONS 0 12330>
 "00000000000000000011000000101011", -- 12330 FREE #<CONS 0 12331>
 "00000000000000000011000000101100", -- 12331 FREE #<CONS 0 12332>
 "00000000000000000011000000101101", -- 12332 FREE #<CONS 0 12333>
 "00000000000000000011000000101110", -- 12333 FREE #<CONS 0 12334>
 "00000000000000000011000000101111", -- 12334 FREE #<CONS 0 12335>
 "00000000000000000011000000110000", -- 12335 FREE #<CONS 0 12336>
 "00000000000000000011000000110001", -- 12336 FREE #<CONS 0 12337>
 "00000000000000000011000000110010", -- 12337 FREE #<CONS 0 12338>
 "00000000000000000011000000110011", -- 12338 FREE #<CONS 0 12339>
 "00000000000000000011000000110100", -- 12339 FREE #<CONS 0 12340>
 "00000000000000000011000000110101", -- 12340 FREE #<CONS 0 12341>
 "00000000000000000011000000110110", -- 12341 FREE #<CONS 0 12342>
 "00000000000000000011000000110111", -- 12342 FREE #<CONS 0 12343>
 "00000000000000000011000000111000", -- 12343 FREE #<CONS 0 12344>
 "00000000000000000011000000111001", -- 12344 FREE #<CONS 0 12345>
 "00000000000000000011000000111010", -- 12345 FREE #<CONS 0 12346>
 "00000000000000000011000000111011", -- 12346 FREE #<CONS 0 12347>
 "00000000000000000011000000111100", -- 12347 FREE #<CONS 0 12348>
 "00000000000000000011000000111101", -- 12348 FREE #<CONS 0 12349>
 "00000000000000000011000000111110", -- 12349 FREE #<CONS 0 12350>
 "00000000000000000011000000111111", -- 12350 FREE #<CONS 0 12351>
 "00000000000000000011000001000000", -- 12351 FREE #<CONS 0 12352>
 "00000000000000000011000001000001", -- 12352 FREE #<CONS 0 12353>
 "00000000000000000011000001000010", -- 12353 FREE #<CONS 0 12354>
 "00000000000000000011000001000011", -- 12354 FREE #<CONS 0 12355>
 "00000000000000000011000001000100", -- 12355 FREE #<CONS 0 12356>
 "00000000000000000011000001000101", -- 12356 FREE #<CONS 0 12357>
 "00000000000000000011000001000110", -- 12357 FREE #<CONS 0 12358>
 "00000000000000000011000001000111", -- 12358 FREE #<CONS 0 12359>
 "00000000000000000011000001001000", -- 12359 FREE #<CONS 0 12360>
 "00000000000000000011000001001001", -- 12360 FREE #<CONS 0 12361>
 "00000000000000000011000001001010", -- 12361 FREE #<CONS 0 12362>
 "00000000000000000011000001001011", -- 12362 FREE #<CONS 0 12363>
 "00000000000000000011000001001100", -- 12363 FREE #<CONS 0 12364>
 "00000000000000000011000001001101", -- 12364 FREE #<CONS 0 12365>
 "00000000000000000011000001001110", -- 12365 FREE #<CONS 0 12366>
 "00000000000000000011000001001111", -- 12366 FREE #<CONS 0 12367>
 "00000000000000000011000001010000", -- 12367 FREE #<CONS 0 12368>
 "00000000000000000011000001010001", -- 12368 FREE #<CONS 0 12369>
 "00000000000000000011000001010010", -- 12369 FREE #<CONS 0 12370>
 "00000000000000000011000001010011", -- 12370 FREE #<CONS 0 12371>
 "00000000000000000011000001010100", -- 12371 FREE #<CONS 0 12372>
 "00000000000000000011000001010101", -- 12372 FREE #<CONS 0 12373>
 "00000000000000000011000001010110", -- 12373 FREE #<CONS 0 12374>
 "00000000000000000011000001010111", -- 12374 FREE #<CONS 0 12375>
 "00000000000000000011000001011000", -- 12375 FREE #<CONS 0 12376>
 "00000000000000000011000001011001", -- 12376 FREE #<CONS 0 12377>
 "00000000000000000011000001011010", -- 12377 FREE #<CONS 0 12378>
 "00000000000000000011000001011011", -- 12378 FREE #<CONS 0 12379>
 "00000000000000000011000001011100", -- 12379 FREE #<CONS 0 12380>
 "00000000000000000011000001011101", -- 12380 FREE #<CONS 0 12381>
 "00000000000000000011000001011110", -- 12381 FREE #<CONS 0 12382>
 "00000000000000000011000001011111", -- 12382 FREE #<CONS 0 12383>
 "00000000000000000011000001100000", -- 12383 FREE #<CONS 0 12384>
 "00000000000000000011000001100001", -- 12384 FREE #<CONS 0 12385>
 "00000000000000000011000001100010", -- 12385 FREE #<CONS 0 12386>
 "00000000000000000011000001100011", -- 12386 FREE #<CONS 0 12387>
 "00000000000000000011000001100100", -- 12387 FREE #<CONS 0 12388>
 "00000000000000000011000001100101", -- 12388 FREE #<CONS 0 12389>
 "00000000000000000011000001100110", -- 12389 FREE #<CONS 0 12390>
 "00000000000000000011000001100111", -- 12390 FREE #<CONS 0 12391>
 "00000000000000000011000001101000", -- 12391 FREE #<CONS 0 12392>
 "00000000000000000011000001101001", -- 12392 FREE #<CONS 0 12393>
 "00000000000000000011000001101010", -- 12393 FREE #<CONS 0 12394>
 "00000000000000000011000001101011", -- 12394 FREE #<CONS 0 12395>
 "00000000000000000011000001101100", -- 12395 FREE #<CONS 0 12396>
 "00000000000000000011000001101101", -- 12396 FREE #<CONS 0 12397>
 "00000000000000000011000001101110", -- 12397 FREE #<CONS 0 12398>
 "00000000000000000011000001101111", -- 12398 FREE #<CONS 0 12399>
 "00000000000000000011000001110000", -- 12399 FREE #<CONS 0 12400>
 "00000000000000000011000001110001", -- 12400 FREE #<CONS 0 12401>
 "00000000000000000011000001110010", -- 12401 FREE #<CONS 0 12402>
 "00000000000000000011000001110011", -- 12402 FREE #<CONS 0 12403>
 "00000000000000000011000001110100", -- 12403 FREE #<CONS 0 12404>
 "00000000000000000011000001110101", -- 12404 FREE #<CONS 0 12405>
 "00000000000000000011000001110110", -- 12405 FREE #<CONS 0 12406>
 "00000000000000000011000001110111", -- 12406 FREE #<CONS 0 12407>
 "00000000000000000011000001111000", -- 12407 FREE #<CONS 0 12408>
 "00000000000000000011000001111001", -- 12408 FREE #<CONS 0 12409>
 "00000000000000000011000001111010", -- 12409 FREE #<CONS 0 12410>
 "00000000000000000011000001111011", -- 12410 FREE #<CONS 0 12411>
 "00000000000000000011000001111100", -- 12411 FREE #<CONS 0 12412>
 "00000000000000000011000001111101", -- 12412 FREE #<CONS 0 12413>
 "00000000000000000011000001111110", -- 12413 FREE #<CONS 0 12414>
 "00000000000000000011000001111111", -- 12414 FREE #<CONS 0 12415>
 "00000000000000000011000010000000", -- 12415 FREE #<CONS 0 12416>
 "00000000000000000011000010000001", -- 12416 FREE #<CONS 0 12417>
 "00000000000000000011000010000010", -- 12417 FREE #<CONS 0 12418>
 "00000000000000000011000010000011", -- 12418 FREE #<CONS 0 12419>
 "00000000000000000011000010000100", -- 12419 FREE #<CONS 0 12420>
 "00000000000000000011000010000101", -- 12420 FREE #<CONS 0 12421>
 "00000000000000000011000010000110", -- 12421 FREE #<CONS 0 12422>
 "00000000000000000011000010000111", -- 12422 FREE #<CONS 0 12423>
 "00000000000000000011000010001000", -- 12423 FREE #<CONS 0 12424>
 "00000000000000000011000010001001", -- 12424 FREE #<CONS 0 12425>
 "00000000000000000011000010001010", -- 12425 FREE #<CONS 0 12426>
 "00000000000000000011000010001011", -- 12426 FREE #<CONS 0 12427>
 "00000000000000000011000010001100", -- 12427 FREE #<CONS 0 12428>
 "00000000000000000011000010001101", -- 12428 FREE #<CONS 0 12429>
 "00000000000000000011000010001110", -- 12429 FREE #<CONS 0 12430>
 "00000000000000000011000010001111", -- 12430 FREE #<CONS 0 12431>
 "00000000000000000011000010010000", -- 12431 FREE #<CONS 0 12432>
 "00000000000000000011000010010001", -- 12432 FREE #<CONS 0 12433>
 "00000000000000000011000010010010", -- 12433 FREE #<CONS 0 12434>
 "00000000000000000011000010010011", -- 12434 FREE #<CONS 0 12435>
 "00000000000000000011000010010100", -- 12435 FREE #<CONS 0 12436>
 "00000000000000000011000010010101", -- 12436 FREE #<CONS 0 12437>
 "00000000000000000011000010010110", -- 12437 FREE #<CONS 0 12438>
 "00000000000000000011000010010111", -- 12438 FREE #<CONS 0 12439>
 "00000000000000000011000010011000", -- 12439 FREE #<CONS 0 12440>
 "00000000000000000011000010011001", -- 12440 FREE #<CONS 0 12441>
 "00000000000000000011000010011010", -- 12441 FREE #<CONS 0 12442>
 "00000000000000000011000010011011", -- 12442 FREE #<CONS 0 12443>
 "00000000000000000011000010011100", -- 12443 FREE #<CONS 0 12444>
 "00000000000000000011000010011101", -- 12444 FREE #<CONS 0 12445>
 "00000000000000000011000010011110", -- 12445 FREE #<CONS 0 12446>
 "00000000000000000011000010011111", -- 12446 FREE #<CONS 0 12447>
 "00000000000000000011000010100000", -- 12447 FREE #<CONS 0 12448>
 "00000000000000000011000010100001", -- 12448 FREE #<CONS 0 12449>
 "00000000000000000011000010100010", -- 12449 FREE #<CONS 0 12450>
 "00000000000000000011000010100011", -- 12450 FREE #<CONS 0 12451>
 "00000000000000000011000010100100", -- 12451 FREE #<CONS 0 12452>
 "00000000000000000011000010100101", -- 12452 FREE #<CONS 0 12453>
 "00000000000000000011000010100110", -- 12453 FREE #<CONS 0 12454>
 "00000000000000000011000010100111", -- 12454 FREE #<CONS 0 12455>
 "00000000000000000011000010101000", -- 12455 FREE #<CONS 0 12456>
 "00000000000000000011000010101001", -- 12456 FREE #<CONS 0 12457>
 "00000000000000000011000010101010", -- 12457 FREE #<CONS 0 12458>
 "00000000000000000011000010101011", -- 12458 FREE #<CONS 0 12459>
 "00000000000000000011000010101100", -- 12459 FREE #<CONS 0 12460>
 "00000000000000000011000010101101", -- 12460 FREE #<CONS 0 12461>
 "00000000000000000011000010101110", -- 12461 FREE #<CONS 0 12462>
 "00000000000000000011000010101111", -- 12462 FREE #<CONS 0 12463>
 "00000000000000000011000010110000", -- 12463 FREE #<CONS 0 12464>
 "00000000000000000011000010110001", -- 12464 FREE #<CONS 0 12465>
 "00000000000000000011000010110010", -- 12465 FREE #<CONS 0 12466>
 "00000000000000000011000010110011", -- 12466 FREE #<CONS 0 12467>
 "00000000000000000011000010110100", -- 12467 FREE #<CONS 0 12468>
 "00000000000000000011000010110101", -- 12468 FREE #<CONS 0 12469>
 "00000000000000000011000010110110", -- 12469 FREE #<CONS 0 12470>
 "00000000000000000011000010110111", -- 12470 FREE #<CONS 0 12471>
 "00000000000000000011000010111000", -- 12471 FREE #<CONS 0 12472>
 "00000000000000000011000010111001", -- 12472 FREE #<CONS 0 12473>
 "00000000000000000011000010111010", -- 12473 FREE #<CONS 0 12474>
 "00000000000000000011000010111011", -- 12474 FREE #<CONS 0 12475>
 "00000000000000000011000010111100", -- 12475 FREE #<CONS 0 12476>
 "00000000000000000011000010111101", -- 12476 FREE #<CONS 0 12477>
 "00000000000000000011000010111110", -- 12477 FREE #<CONS 0 12478>
 "00000000000000000011000010111111", -- 12478 FREE #<CONS 0 12479>
 "00000000000000000011000011000000", -- 12479 FREE #<CONS 0 12480>
 "00000000000000000011000011000001", -- 12480 FREE #<CONS 0 12481>
 "00000000000000000011000011000010", -- 12481 FREE #<CONS 0 12482>
 "00000000000000000011000011000011", -- 12482 FREE #<CONS 0 12483>
 "00000000000000000011000011000100", -- 12483 FREE #<CONS 0 12484>
 "00000000000000000011000011000101", -- 12484 FREE #<CONS 0 12485>
 "00000000000000000011000011000110", -- 12485 FREE #<CONS 0 12486>
 "00000000000000000011000011000111", -- 12486 FREE #<CONS 0 12487>
 "00000000000000000011000011001000", -- 12487 FREE #<CONS 0 12488>
 "00000000000000000011000011001001", -- 12488 FREE #<CONS 0 12489>
 "00000000000000000011000011001010", -- 12489 FREE #<CONS 0 12490>
 "00000000000000000011000011001011", -- 12490 FREE #<CONS 0 12491>
 "00000000000000000011000011001100", -- 12491 FREE #<CONS 0 12492>
 "00000000000000000011000011001101", -- 12492 FREE #<CONS 0 12493>
 "00000000000000000011000011001110", -- 12493 FREE #<CONS 0 12494>
 "00000000000000000011000011001111", -- 12494 FREE #<CONS 0 12495>
 "00000000000000000011000011010000", -- 12495 FREE #<CONS 0 12496>
 "00000000000000000011000011010001", -- 12496 FREE #<CONS 0 12497>
 "00000000000000000011000011010010", -- 12497 FREE #<CONS 0 12498>
 "00000000000000000011000011010011", -- 12498 FREE #<CONS 0 12499>
 "00000000000000000011000011010100", -- 12499 FREE #<CONS 0 12500>
 "00000000000000000011000011010101", -- 12500 FREE #<CONS 0 12501>
 "00000000000000000011000011010110", -- 12501 FREE #<CONS 0 12502>
 "00000000000000000011000011010111", -- 12502 FREE #<CONS 0 12503>
 "00000000000000000011000011011000", -- 12503 FREE #<CONS 0 12504>
 "00000000000000000011000011011001", -- 12504 FREE #<CONS 0 12505>
 "00000000000000000011000011011010", -- 12505 FREE #<CONS 0 12506>
 "00000000000000000011000011011011", -- 12506 FREE #<CONS 0 12507>
 "00000000000000000011000011011100", -- 12507 FREE #<CONS 0 12508>
 "00000000000000000011000011011101", -- 12508 FREE #<CONS 0 12509>
 "00000000000000000011000011011110", -- 12509 FREE #<CONS 0 12510>
 "00000000000000000011000011011111", -- 12510 FREE #<CONS 0 12511>
 "00000000000000000011000011100000", -- 12511 FREE #<CONS 0 12512>
 "00000000000000000011000011100001", -- 12512 FREE #<CONS 0 12513>
 "00000000000000000011000011100010", -- 12513 FREE #<CONS 0 12514>
 "00000000000000000011000011100011", -- 12514 FREE #<CONS 0 12515>
 "00000000000000000011000011100100", -- 12515 FREE #<CONS 0 12516>
 "00000000000000000011000011100101", -- 12516 FREE #<CONS 0 12517>
 "00000000000000000011000011100110", -- 12517 FREE #<CONS 0 12518>
 "00000000000000000011000011100111", -- 12518 FREE #<CONS 0 12519>
 "00000000000000000011000011101000", -- 12519 FREE #<CONS 0 12520>
 "00000000000000000011000011101001", -- 12520 FREE #<CONS 0 12521>
 "00000000000000000011000011101010", -- 12521 FREE #<CONS 0 12522>
 "00000000000000000011000011101011", -- 12522 FREE #<CONS 0 12523>
 "00000000000000000011000011101100", -- 12523 FREE #<CONS 0 12524>
 "00000000000000000011000011101101", -- 12524 FREE #<CONS 0 12525>
 "00000000000000000011000011101110", -- 12525 FREE #<CONS 0 12526>
 "00000000000000000011000011101111", -- 12526 FREE #<CONS 0 12527>
 "00000000000000000011000011110000", -- 12527 FREE #<CONS 0 12528>
 "00000000000000000011000011110001", -- 12528 FREE #<CONS 0 12529>
 "00000000000000000011000011110010", -- 12529 FREE #<CONS 0 12530>
 "00000000000000000011000011110011", -- 12530 FREE #<CONS 0 12531>
 "00000000000000000011000011110100", -- 12531 FREE #<CONS 0 12532>
 "00000000000000000011000011110101", -- 12532 FREE #<CONS 0 12533>
 "00000000000000000011000011110110", -- 12533 FREE #<CONS 0 12534>
 "00000000000000000011000011110111", -- 12534 FREE #<CONS 0 12535>
 "00000000000000000011000011111000", -- 12535 FREE #<CONS 0 12536>
 "00000000000000000011000011111001", -- 12536 FREE #<CONS 0 12537>
 "00000000000000000011000011111010", -- 12537 FREE #<CONS 0 12538>
 "00000000000000000011000011111011", -- 12538 FREE #<CONS 0 12539>
 "00000000000000000011000011111100", -- 12539 FREE #<CONS 0 12540>
 "00000000000000000011000011111101", -- 12540 FREE #<CONS 0 12541>
 "00000000000000000011000011111110", -- 12541 FREE #<CONS 0 12542>
 "00000000000000000011000011111111", -- 12542 FREE #<CONS 0 12543>
 "00000000000000000011000100000000", -- 12543 FREE #<CONS 0 12544>
 "00000000000000000011000100000001", -- 12544 FREE #<CONS 0 12545>
 "00000000000000000011000100000010", -- 12545 FREE #<CONS 0 12546>
 "00000000000000000011000100000011", -- 12546 FREE #<CONS 0 12547>
 "00000000000000000011000100000100", -- 12547 FREE #<CONS 0 12548>
 "00000000000000000011000100000101", -- 12548 FREE #<CONS 0 12549>
 "00000000000000000011000100000110", -- 12549 FREE #<CONS 0 12550>
 "00000000000000000011000100000111", -- 12550 FREE #<CONS 0 12551>
 "00000000000000000011000100001000", -- 12551 FREE #<CONS 0 12552>
 "00000000000000000011000100001001", -- 12552 FREE #<CONS 0 12553>
 "00000000000000000011000100001010", -- 12553 FREE #<CONS 0 12554>
 "00000000000000000011000100001011", -- 12554 FREE #<CONS 0 12555>
 "00000000000000000011000100001100", -- 12555 FREE #<CONS 0 12556>
 "00000000000000000011000100001101", -- 12556 FREE #<CONS 0 12557>
 "00000000000000000011000100001110", -- 12557 FREE #<CONS 0 12558>
 "00000000000000000011000100001111", -- 12558 FREE #<CONS 0 12559>
 "00000000000000000011000100010000", -- 12559 FREE #<CONS 0 12560>
 "00000000000000000011000100010001", -- 12560 FREE #<CONS 0 12561>
 "00000000000000000011000100010010", -- 12561 FREE #<CONS 0 12562>
 "00000000000000000011000100010011", -- 12562 FREE #<CONS 0 12563>
 "00000000000000000011000100010100", -- 12563 FREE #<CONS 0 12564>
 "00000000000000000011000100010101", -- 12564 FREE #<CONS 0 12565>
 "00000000000000000011000100010110", -- 12565 FREE #<CONS 0 12566>
 "00000000000000000011000100010111", -- 12566 FREE #<CONS 0 12567>
 "00000000000000000011000100011000", -- 12567 FREE #<CONS 0 12568>
 "00000000000000000011000100011001", -- 12568 FREE #<CONS 0 12569>
 "00000000000000000011000100011010", -- 12569 FREE #<CONS 0 12570>
 "00000000000000000011000100011011", -- 12570 FREE #<CONS 0 12571>
 "00000000000000000011000100011100", -- 12571 FREE #<CONS 0 12572>
 "00000000000000000011000100011101", -- 12572 FREE #<CONS 0 12573>
 "00000000000000000011000100011110", -- 12573 FREE #<CONS 0 12574>
 "00000000000000000011000100011111", -- 12574 FREE #<CONS 0 12575>
 "00000000000000000011000100100000", -- 12575 FREE #<CONS 0 12576>
 "00000000000000000011000100100001", -- 12576 FREE #<CONS 0 12577>
 "00000000000000000011000100100010", -- 12577 FREE #<CONS 0 12578>
 "00000000000000000011000100100011", -- 12578 FREE #<CONS 0 12579>
 "00000000000000000011000100100100", -- 12579 FREE #<CONS 0 12580>
 "00000000000000000011000100100101", -- 12580 FREE #<CONS 0 12581>
 "00000000000000000011000100100110", -- 12581 FREE #<CONS 0 12582>
 "00000000000000000011000100100111", -- 12582 FREE #<CONS 0 12583>
 "00000000000000000011000100101000", -- 12583 FREE #<CONS 0 12584>
 "00000000000000000011000100101001", -- 12584 FREE #<CONS 0 12585>
 "00000000000000000011000100101010", -- 12585 FREE #<CONS 0 12586>
 "00000000000000000011000100101011", -- 12586 FREE #<CONS 0 12587>
 "00000000000000000011000100101100", -- 12587 FREE #<CONS 0 12588>
 "00000000000000000011000100101101", -- 12588 FREE #<CONS 0 12589>
 "00000000000000000011000100101110", -- 12589 FREE #<CONS 0 12590>
 "00000000000000000011000100101111", -- 12590 FREE #<CONS 0 12591>
 "00000000000000000011000100110000", -- 12591 FREE #<CONS 0 12592>
 "00000000000000000011000100110001", -- 12592 FREE #<CONS 0 12593>
 "00000000000000000011000100110010", -- 12593 FREE #<CONS 0 12594>
 "00000000000000000011000100110011", -- 12594 FREE #<CONS 0 12595>
 "00000000000000000011000100110100", -- 12595 FREE #<CONS 0 12596>
 "00000000000000000011000100110101", -- 12596 FREE #<CONS 0 12597>
 "00000000000000000011000100110110", -- 12597 FREE #<CONS 0 12598>
 "00000000000000000011000100110111", -- 12598 FREE #<CONS 0 12599>
 "00000000000000000011000100111000", -- 12599 FREE #<CONS 0 12600>
 "00000000000000000011000100111001", -- 12600 FREE #<CONS 0 12601>
 "00000000000000000011000100111010", -- 12601 FREE #<CONS 0 12602>
 "00000000000000000011000100111011", -- 12602 FREE #<CONS 0 12603>
 "00000000000000000011000100111100", -- 12603 FREE #<CONS 0 12604>
 "00000000000000000011000100111101", -- 12604 FREE #<CONS 0 12605>
 "00000000000000000011000100111110", -- 12605 FREE #<CONS 0 12606>
 "00000000000000000011000100111111", -- 12606 FREE #<CONS 0 12607>
 "00000000000000000011000101000000", -- 12607 FREE #<CONS 0 12608>
 "00000000000000000011000101000001", -- 12608 FREE #<CONS 0 12609>
 "00000000000000000011000101000010", -- 12609 FREE #<CONS 0 12610>
 "00000000000000000011000101000011", -- 12610 FREE #<CONS 0 12611>
 "00000000000000000011000101000100", -- 12611 FREE #<CONS 0 12612>
 "00000000000000000011000101000101", -- 12612 FREE #<CONS 0 12613>
 "00000000000000000011000101000110", -- 12613 FREE #<CONS 0 12614>
 "00000000000000000011000101000111", -- 12614 FREE #<CONS 0 12615>
 "00000000000000000011000101001000", -- 12615 FREE #<CONS 0 12616>
 "00000000000000000011000101001001", -- 12616 FREE #<CONS 0 12617>
 "00000000000000000011000101001010", -- 12617 FREE #<CONS 0 12618>
 "00000000000000000011000101001011", -- 12618 FREE #<CONS 0 12619>
 "00000000000000000011000101001100", -- 12619 FREE #<CONS 0 12620>
 "00000000000000000011000101001101", -- 12620 FREE #<CONS 0 12621>
 "00000000000000000011000101001110", -- 12621 FREE #<CONS 0 12622>
 "00000000000000000011000101001111", -- 12622 FREE #<CONS 0 12623>
 "00000000000000000011000101010000", -- 12623 FREE #<CONS 0 12624>
 "00000000000000000011000101010001", -- 12624 FREE #<CONS 0 12625>
 "00000000000000000011000101010010", -- 12625 FREE #<CONS 0 12626>
 "00000000000000000011000101010011", -- 12626 FREE #<CONS 0 12627>
 "00000000000000000011000101010100", -- 12627 FREE #<CONS 0 12628>
 "00000000000000000011000101010101", -- 12628 FREE #<CONS 0 12629>
 "00000000000000000011000101010110", -- 12629 FREE #<CONS 0 12630>
 "00000000000000000011000101010111", -- 12630 FREE #<CONS 0 12631>
 "00000000000000000011000101011000", -- 12631 FREE #<CONS 0 12632>
 "00000000000000000011000101011001", -- 12632 FREE #<CONS 0 12633>
 "00000000000000000011000101011010", -- 12633 FREE #<CONS 0 12634>
 "00000000000000000011000101011011", -- 12634 FREE #<CONS 0 12635>
 "00000000000000000011000101011100", -- 12635 FREE #<CONS 0 12636>
 "00000000000000000011000101011101", -- 12636 FREE #<CONS 0 12637>
 "00000000000000000011000101011110", -- 12637 FREE #<CONS 0 12638>
 "00000000000000000011000101011111", -- 12638 FREE #<CONS 0 12639>
 "00000000000000000011000101100000", -- 12639 FREE #<CONS 0 12640>
 "00000000000000000011000101100001", -- 12640 FREE #<CONS 0 12641>
 "00000000000000000011000101100010", -- 12641 FREE #<CONS 0 12642>
 "00000000000000000011000101100011", -- 12642 FREE #<CONS 0 12643>
 "00000000000000000011000101100100", -- 12643 FREE #<CONS 0 12644>
 "00000000000000000011000101100101", -- 12644 FREE #<CONS 0 12645>
 "00000000000000000011000101100110", -- 12645 FREE #<CONS 0 12646>
 "00000000000000000011000101100111", -- 12646 FREE #<CONS 0 12647>
 "00000000000000000011000101101000", -- 12647 FREE #<CONS 0 12648>
 "00000000000000000011000101101001", -- 12648 FREE #<CONS 0 12649>
 "00000000000000000011000101101010", -- 12649 FREE #<CONS 0 12650>
 "00000000000000000011000101101011", -- 12650 FREE #<CONS 0 12651>
 "00000000000000000011000101101100", -- 12651 FREE #<CONS 0 12652>
 "00000000000000000011000101101101", -- 12652 FREE #<CONS 0 12653>
 "00000000000000000011000101101110", -- 12653 FREE #<CONS 0 12654>
 "00000000000000000011000101101111", -- 12654 FREE #<CONS 0 12655>
 "00000000000000000011000101110000", -- 12655 FREE #<CONS 0 12656>
 "00000000000000000011000101110001", -- 12656 FREE #<CONS 0 12657>
 "00000000000000000011000101110010", -- 12657 FREE #<CONS 0 12658>
 "00000000000000000011000101110011", -- 12658 FREE #<CONS 0 12659>
 "00000000000000000011000101110100", -- 12659 FREE #<CONS 0 12660>
 "00000000000000000011000101110101", -- 12660 FREE #<CONS 0 12661>
 "00000000000000000011000101110110", -- 12661 FREE #<CONS 0 12662>
 "00000000000000000011000101110111", -- 12662 FREE #<CONS 0 12663>
 "00000000000000000011000101111000", -- 12663 FREE #<CONS 0 12664>
 "00000000000000000011000101111001", -- 12664 FREE #<CONS 0 12665>
 "00000000000000000011000101111010", -- 12665 FREE #<CONS 0 12666>
 "00000000000000000011000101111011", -- 12666 FREE #<CONS 0 12667>
 "00000000000000000011000101111100", -- 12667 FREE #<CONS 0 12668>
 "00000000000000000011000101111101", -- 12668 FREE #<CONS 0 12669>
 "00000000000000000011000101111110", -- 12669 FREE #<CONS 0 12670>
 "00000000000000000011000101111111", -- 12670 FREE #<CONS 0 12671>
 "00000000000000000011000110000000", -- 12671 FREE #<CONS 0 12672>
 "00000000000000000011000110000001", -- 12672 FREE #<CONS 0 12673>
 "00000000000000000011000110000010", -- 12673 FREE #<CONS 0 12674>
 "00000000000000000011000110000011", -- 12674 FREE #<CONS 0 12675>
 "00000000000000000011000110000100", -- 12675 FREE #<CONS 0 12676>
 "00000000000000000011000110000101", -- 12676 FREE #<CONS 0 12677>
 "00000000000000000011000110000110", -- 12677 FREE #<CONS 0 12678>
 "00000000000000000011000110000111", -- 12678 FREE #<CONS 0 12679>
 "00000000000000000011000110001000", -- 12679 FREE #<CONS 0 12680>
 "00000000000000000011000110001001", -- 12680 FREE #<CONS 0 12681>
 "00000000000000000011000110001010", -- 12681 FREE #<CONS 0 12682>
 "00000000000000000011000110001011", -- 12682 FREE #<CONS 0 12683>
 "00000000000000000011000110001100", -- 12683 FREE #<CONS 0 12684>
 "00000000000000000011000110001101", -- 12684 FREE #<CONS 0 12685>
 "00000000000000000011000110001110", -- 12685 FREE #<CONS 0 12686>
 "00000000000000000011000110001111", -- 12686 FREE #<CONS 0 12687>
 "00000000000000000011000110010000", -- 12687 FREE #<CONS 0 12688>
 "00000000000000000011000110010001", -- 12688 FREE #<CONS 0 12689>
 "00000000000000000011000110010010", -- 12689 FREE #<CONS 0 12690>
 "00000000000000000011000110010011", -- 12690 FREE #<CONS 0 12691>
 "00000000000000000011000110010100", -- 12691 FREE #<CONS 0 12692>
 "00000000000000000011000110010101", -- 12692 FREE #<CONS 0 12693>
 "00000000000000000011000110010110", -- 12693 FREE #<CONS 0 12694>
 "00000000000000000011000110010111", -- 12694 FREE #<CONS 0 12695>
 "00000000000000000011000110011000", -- 12695 FREE #<CONS 0 12696>
 "00000000000000000011000110011001", -- 12696 FREE #<CONS 0 12697>
 "00000000000000000011000110011010", -- 12697 FREE #<CONS 0 12698>
 "00000000000000000011000110011011", -- 12698 FREE #<CONS 0 12699>
 "00000000000000000011000110011100", -- 12699 FREE #<CONS 0 12700>
 "00000000000000000011000110011101", -- 12700 FREE #<CONS 0 12701>
 "00000000000000000011000110011110", -- 12701 FREE #<CONS 0 12702>
 "00000000000000000011000110011111", -- 12702 FREE #<CONS 0 12703>
 "00000000000000000011000110100000", -- 12703 FREE #<CONS 0 12704>
 "00000000000000000011000110100001", -- 12704 FREE #<CONS 0 12705>
 "00000000000000000011000110100010", -- 12705 FREE #<CONS 0 12706>
 "00000000000000000011000110100011", -- 12706 FREE #<CONS 0 12707>
 "00000000000000000011000110100100", -- 12707 FREE #<CONS 0 12708>
 "00000000000000000011000110100101", -- 12708 FREE #<CONS 0 12709>
 "00000000000000000011000110100110", -- 12709 FREE #<CONS 0 12710>
 "00000000000000000011000110100111", -- 12710 FREE #<CONS 0 12711>
 "00000000000000000011000110101000", -- 12711 FREE #<CONS 0 12712>
 "00000000000000000011000110101001", -- 12712 FREE #<CONS 0 12713>
 "00000000000000000011000110101010", -- 12713 FREE #<CONS 0 12714>
 "00000000000000000011000110101011", -- 12714 FREE #<CONS 0 12715>
 "00000000000000000011000110101100", -- 12715 FREE #<CONS 0 12716>
 "00000000000000000011000110101101", -- 12716 FREE #<CONS 0 12717>
 "00000000000000000011000110101110", -- 12717 FREE #<CONS 0 12718>
 "00000000000000000011000110101111", -- 12718 FREE #<CONS 0 12719>
 "00000000000000000011000110110000", -- 12719 FREE #<CONS 0 12720>
 "00000000000000000011000110110001", -- 12720 FREE #<CONS 0 12721>
 "00000000000000000011000110110010", -- 12721 FREE #<CONS 0 12722>
 "00000000000000000011000110110011", -- 12722 FREE #<CONS 0 12723>
 "00000000000000000011000110110100", -- 12723 FREE #<CONS 0 12724>
 "00000000000000000011000110110101", -- 12724 FREE #<CONS 0 12725>
 "00000000000000000011000110110110", -- 12725 FREE #<CONS 0 12726>
 "00000000000000000011000110110111", -- 12726 FREE #<CONS 0 12727>
 "00000000000000000011000110111000", -- 12727 FREE #<CONS 0 12728>
 "00000000000000000011000110111001", -- 12728 FREE #<CONS 0 12729>
 "00000000000000000011000110111010", -- 12729 FREE #<CONS 0 12730>
 "00000000000000000011000110111011", -- 12730 FREE #<CONS 0 12731>
 "00000000000000000011000110111100", -- 12731 FREE #<CONS 0 12732>
 "00000000000000000011000110111101", -- 12732 FREE #<CONS 0 12733>
 "00000000000000000011000110111110", -- 12733 FREE #<CONS 0 12734>
 "00000000000000000011000110111111", -- 12734 FREE #<CONS 0 12735>
 "00000000000000000011000111000000", -- 12735 FREE #<CONS 0 12736>
 "00000000000000000011000111000001", -- 12736 FREE #<CONS 0 12737>
 "00000000000000000011000111000010", -- 12737 FREE #<CONS 0 12738>
 "00000000000000000011000111000011", -- 12738 FREE #<CONS 0 12739>
 "00000000000000000011000111000100", -- 12739 FREE #<CONS 0 12740>
 "00000000000000000011000111000101", -- 12740 FREE #<CONS 0 12741>
 "00000000000000000011000111000110", -- 12741 FREE #<CONS 0 12742>
 "00000000000000000011000111000111", -- 12742 FREE #<CONS 0 12743>
 "00000000000000000011000111001000", -- 12743 FREE #<CONS 0 12744>
 "00000000000000000011000111001001", -- 12744 FREE #<CONS 0 12745>
 "00000000000000000011000111001010", -- 12745 FREE #<CONS 0 12746>
 "00000000000000000011000111001011", -- 12746 FREE #<CONS 0 12747>
 "00000000000000000011000111001100", -- 12747 FREE #<CONS 0 12748>
 "00000000000000000011000111001101", -- 12748 FREE #<CONS 0 12749>
 "00000000000000000011000111001110", -- 12749 FREE #<CONS 0 12750>
 "00000000000000000011000111001111", -- 12750 FREE #<CONS 0 12751>
 "00000000000000000011000111010000", -- 12751 FREE #<CONS 0 12752>
 "00000000000000000011000111010001", -- 12752 FREE #<CONS 0 12753>
 "00000000000000000011000111010010", -- 12753 FREE #<CONS 0 12754>
 "00000000000000000011000111010011", -- 12754 FREE #<CONS 0 12755>
 "00000000000000000011000111010100", -- 12755 FREE #<CONS 0 12756>
 "00000000000000000011000111010101", -- 12756 FREE #<CONS 0 12757>
 "00000000000000000011000111010110", -- 12757 FREE #<CONS 0 12758>
 "00000000000000000011000111010111", -- 12758 FREE #<CONS 0 12759>
 "00000000000000000011000111011000", -- 12759 FREE #<CONS 0 12760>
 "00000000000000000011000111011001", -- 12760 FREE #<CONS 0 12761>
 "00000000000000000011000111011010", -- 12761 FREE #<CONS 0 12762>
 "00000000000000000011000111011011", -- 12762 FREE #<CONS 0 12763>
 "00000000000000000011000111011100", -- 12763 FREE #<CONS 0 12764>
 "00000000000000000011000111011101", -- 12764 FREE #<CONS 0 12765>
 "00000000000000000011000111011110", -- 12765 FREE #<CONS 0 12766>
 "00000000000000000011000111011111", -- 12766 FREE #<CONS 0 12767>
 "00000000000000000011000111100000", -- 12767 FREE #<CONS 0 12768>
 "00000000000000000011000111100001", -- 12768 FREE #<CONS 0 12769>
 "00000000000000000011000111100010", -- 12769 FREE #<CONS 0 12770>
 "00000000000000000011000111100011", -- 12770 FREE #<CONS 0 12771>
 "00000000000000000011000111100100", -- 12771 FREE #<CONS 0 12772>
 "00000000000000000011000111100101", -- 12772 FREE #<CONS 0 12773>
 "00000000000000000011000111100110", -- 12773 FREE #<CONS 0 12774>
 "00000000000000000011000111100111", -- 12774 FREE #<CONS 0 12775>
 "00000000000000000011000111101000", -- 12775 FREE #<CONS 0 12776>
 "00000000000000000011000111101001", -- 12776 FREE #<CONS 0 12777>
 "00000000000000000011000111101010", -- 12777 FREE #<CONS 0 12778>
 "00000000000000000011000111101011", -- 12778 FREE #<CONS 0 12779>
 "00000000000000000011000111101100", -- 12779 FREE #<CONS 0 12780>
 "00000000000000000011000111101101", -- 12780 FREE #<CONS 0 12781>
 "00000000000000000011000111101110", -- 12781 FREE #<CONS 0 12782>
 "00000000000000000011000111101111", -- 12782 FREE #<CONS 0 12783>
 "00000000000000000011000111110000", -- 12783 FREE #<CONS 0 12784>
 "00000000000000000011000111110001", -- 12784 FREE #<CONS 0 12785>
 "00000000000000000011000111110010", -- 12785 FREE #<CONS 0 12786>
 "00000000000000000011000111110011", -- 12786 FREE #<CONS 0 12787>
 "00000000000000000011000111110100", -- 12787 FREE #<CONS 0 12788>
 "00000000000000000011000111110101", -- 12788 FREE #<CONS 0 12789>
 "00000000000000000011000111110110", -- 12789 FREE #<CONS 0 12790>
 "00000000000000000011000111110111", -- 12790 FREE #<CONS 0 12791>
 "00000000000000000011000111111000", -- 12791 FREE #<CONS 0 12792>
 "00000000000000000011000111111001", -- 12792 FREE #<CONS 0 12793>
 "00000000000000000011000111111010", -- 12793 FREE #<CONS 0 12794>
 "00000000000000000011000111111011", -- 12794 FREE #<CONS 0 12795>
 "00000000000000000011000111111100", -- 12795 FREE #<CONS 0 12796>
 "00000000000000000011000111111101", -- 12796 FREE #<CONS 0 12797>
 "00000000000000000011000111111110", -- 12797 FREE #<CONS 0 12798>
 "00000000000000000011000111111111", -- 12798 FREE #<CONS 0 12799>
 "00000000000000000011001000000000", -- 12799 FREE #<CONS 0 12800>
 "00000000000000000011001000000001", -- 12800 FREE #<CONS 0 12801>
 "00000000000000000011001000000010", -- 12801 FREE #<CONS 0 12802>
 "00000000000000000011001000000011", -- 12802 FREE #<CONS 0 12803>
 "00000000000000000011001000000100", -- 12803 FREE #<CONS 0 12804>
 "00000000000000000011001000000101", -- 12804 FREE #<CONS 0 12805>
 "00000000000000000011001000000110", -- 12805 FREE #<CONS 0 12806>
 "00000000000000000011001000000111", -- 12806 FREE #<CONS 0 12807>
 "00000000000000000011001000001000", -- 12807 FREE #<CONS 0 12808>
 "00000000000000000011001000001001", -- 12808 FREE #<CONS 0 12809>
 "00000000000000000011001000001010", -- 12809 FREE #<CONS 0 12810>
 "00000000000000000011001000001011", -- 12810 FREE #<CONS 0 12811>
 "00000000000000000011001000001100", -- 12811 FREE #<CONS 0 12812>
 "00000000000000000011001000001101", -- 12812 FREE #<CONS 0 12813>
 "00000000000000000011001000001110", -- 12813 FREE #<CONS 0 12814>
 "00000000000000000011001000001111", -- 12814 FREE #<CONS 0 12815>
 "00000000000000000011001000010000", -- 12815 FREE #<CONS 0 12816>
 "00000000000000000011001000010001", -- 12816 FREE #<CONS 0 12817>
 "00000000000000000011001000010010", -- 12817 FREE #<CONS 0 12818>
 "00000000000000000011001000010011", -- 12818 FREE #<CONS 0 12819>
 "00000000000000000011001000010100", -- 12819 FREE #<CONS 0 12820>
 "00000000000000000011001000010101", -- 12820 FREE #<CONS 0 12821>
 "00000000000000000011001000010110", -- 12821 FREE #<CONS 0 12822>
 "00000000000000000011001000010111", -- 12822 FREE #<CONS 0 12823>
 "00000000000000000011001000011000", -- 12823 FREE #<CONS 0 12824>
 "00000000000000000011001000011001", -- 12824 FREE #<CONS 0 12825>
 "00000000000000000011001000011010", -- 12825 FREE #<CONS 0 12826>
 "00000000000000000011001000011011", -- 12826 FREE #<CONS 0 12827>
 "00000000000000000011001000011100", -- 12827 FREE #<CONS 0 12828>
 "00000000000000000011001000011101", -- 12828 FREE #<CONS 0 12829>
 "00000000000000000011001000011110", -- 12829 FREE #<CONS 0 12830>
 "00000000000000000011001000011111", -- 12830 FREE #<CONS 0 12831>
 "00000000000000000011001000100000", -- 12831 FREE #<CONS 0 12832>
 "00000000000000000011001000100001", -- 12832 FREE #<CONS 0 12833>
 "00000000000000000011001000100010", -- 12833 FREE #<CONS 0 12834>
 "00000000000000000011001000100011", -- 12834 FREE #<CONS 0 12835>
 "00000000000000000011001000100100", -- 12835 FREE #<CONS 0 12836>
 "00000000000000000011001000100101", -- 12836 FREE #<CONS 0 12837>
 "00000000000000000011001000100110", -- 12837 FREE #<CONS 0 12838>
 "00000000000000000011001000100111", -- 12838 FREE #<CONS 0 12839>
 "00000000000000000011001000101000", -- 12839 FREE #<CONS 0 12840>
 "00000000000000000011001000101001", -- 12840 FREE #<CONS 0 12841>
 "00000000000000000011001000101010", -- 12841 FREE #<CONS 0 12842>
 "00000000000000000011001000101011", -- 12842 FREE #<CONS 0 12843>
 "00000000000000000011001000101100", -- 12843 FREE #<CONS 0 12844>
 "00000000000000000011001000101101", -- 12844 FREE #<CONS 0 12845>
 "00000000000000000011001000101110", -- 12845 FREE #<CONS 0 12846>
 "00000000000000000011001000101111", -- 12846 FREE #<CONS 0 12847>
 "00000000000000000011001000110000", -- 12847 FREE #<CONS 0 12848>
 "00000000000000000011001000110001", -- 12848 FREE #<CONS 0 12849>
 "00000000000000000011001000110010", -- 12849 FREE #<CONS 0 12850>
 "00000000000000000011001000110011", -- 12850 FREE #<CONS 0 12851>
 "00000000000000000011001000110100", -- 12851 FREE #<CONS 0 12852>
 "00000000000000000011001000110101", -- 12852 FREE #<CONS 0 12853>
 "00000000000000000011001000110110", -- 12853 FREE #<CONS 0 12854>
 "00000000000000000011001000110111", -- 12854 FREE #<CONS 0 12855>
 "00000000000000000011001000111000", -- 12855 FREE #<CONS 0 12856>
 "00000000000000000011001000111001", -- 12856 FREE #<CONS 0 12857>
 "00000000000000000011001000111010", -- 12857 FREE #<CONS 0 12858>
 "00000000000000000011001000111011", -- 12858 FREE #<CONS 0 12859>
 "00000000000000000011001000111100", -- 12859 FREE #<CONS 0 12860>
 "00000000000000000011001000111101", -- 12860 FREE #<CONS 0 12861>
 "00000000000000000011001000111110", -- 12861 FREE #<CONS 0 12862>
 "00000000000000000011001000111111", -- 12862 FREE #<CONS 0 12863>
 "00000000000000000011001001000000", -- 12863 FREE #<CONS 0 12864>
 "00000000000000000011001001000001", -- 12864 FREE #<CONS 0 12865>
 "00000000000000000011001001000010", -- 12865 FREE #<CONS 0 12866>
 "00000000000000000011001001000011", -- 12866 FREE #<CONS 0 12867>
 "00000000000000000011001001000100", -- 12867 FREE #<CONS 0 12868>
 "00000000000000000011001001000101", -- 12868 FREE #<CONS 0 12869>
 "00000000000000000011001001000110", -- 12869 FREE #<CONS 0 12870>
 "00000000000000000011001001000111", -- 12870 FREE #<CONS 0 12871>
 "00000000000000000011001001001000", -- 12871 FREE #<CONS 0 12872>
 "00000000000000000011001001001001", -- 12872 FREE #<CONS 0 12873>
 "00000000000000000011001001001010", -- 12873 FREE #<CONS 0 12874>
 "00000000000000000011001001001011", -- 12874 FREE #<CONS 0 12875>
 "00000000000000000011001001001100", -- 12875 FREE #<CONS 0 12876>
 "00000000000000000011001001001101", -- 12876 FREE #<CONS 0 12877>
 "00000000000000000011001001001110", -- 12877 FREE #<CONS 0 12878>
 "00000000000000000011001001001111", -- 12878 FREE #<CONS 0 12879>
 "00000000000000000011001001010000", -- 12879 FREE #<CONS 0 12880>
 "00000000000000000011001001010001", -- 12880 FREE #<CONS 0 12881>
 "00000000000000000011001001010010", -- 12881 FREE #<CONS 0 12882>
 "00000000000000000011001001010011", -- 12882 FREE #<CONS 0 12883>
 "00000000000000000011001001010100", -- 12883 FREE #<CONS 0 12884>
 "00000000000000000011001001010101", -- 12884 FREE #<CONS 0 12885>
 "00000000000000000011001001010110", -- 12885 FREE #<CONS 0 12886>
 "00000000000000000011001001010111", -- 12886 FREE #<CONS 0 12887>
 "00000000000000000011001001011000", -- 12887 FREE #<CONS 0 12888>
 "00000000000000000011001001011001", -- 12888 FREE #<CONS 0 12889>
 "00000000000000000011001001011010", -- 12889 FREE #<CONS 0 12890>
 "00000000000000000011001001011011", -- 12890 FREE #<CONS 0 12891>
 "00000000000000000011001001011100", -- 12891 FREE #<CONS 0 12892>
 "00000000000000000011001001011101", -- 12892 FREE #<CONS 0 12893>
 "00000000000000000011001001011110", -- 12893 FREE #<CONS 0 12894>
 "00000000000000000011001001011111", -- 12894 FREE #<CONS 0 12895>
 "00000000000000000011001001100000", -- 12895 FREE #<CONS 0 12896>
 "00000000000000000011001001100001", -- 12896 FREE #<CONS 0 12897>
 "00000000000000000011001001100010", -- 12897 FREE #<CONS 0 12898>
 "00000000000000000011001001100011", -- 12898 FREE #<CONS 0 12899>
 "00000000000000000011001001100100", -- 12899 FREE #<CONS 0 12900>
 "00000000000000000011001001100101", -- 12900 FREE #<CONS 0 12901>
 "00000000000000000011001001100110", -- 12901 FREE #<CONS 0 12902>
 "00000000000000000011001001100111", -- 12902 FREE #<CONS 0 12903>
 "00000000000000000011001001101000", -- 12903 FREE #<CONS 0 12904>
 "00000000000000000011001001101001", -- 12904 FREE #<CONS 0 12905>
 "00000000000000000011001001101010", -- 12905 FREE #<CONS 0 12906>
 "00000000000000000011001001101011", -- 12906 FREE #<CONS 0 12907>
 "00000000000000000011001001101100", -- 12907 FREE #<CONS 0 12908>
 "00000000000000000011001001101101", -- 12908 FREE #<CONS 0 12909>
 "00000000000000000011001001101110", -- 12909 FREE #<CONS 0 12910>
 "00000000000000000011001001101111", -- 12910 FREE #<CONS 0 12911>
 "00000000000000000011001001110000", -- 12911 FREE #<CONS 0 12912>
 "00000000000000000011001001110001", -- 12912 FREE #<CONS 0 12913>
 "00000000000000000011001001110010", -- 12913 FREE #<CONS 0 12914>
 "00000000000000000011001001110011", -- 12914 FREE #<CONS 0 12915>
 "00000000000000000011001001110100", -- 12915 FREE #<CONS 0 12916>
 "00000000000000000011001001110101", -- 12916 FREE #<CONS 0 12917>
 "00000000000000000011001001110110", -- 12917 FREE #<CONS 0 12918>
 "00000000000000000011001001110111", -- 12918 FREE #<CONS 0 12919>
 "00000000000000000011001001111000", -- 12919 FREE #<CONS 0 12920>
 "00000000000000000011001001111001", -- 12920 FREE #<CONS 0 12921>
 "00000000000000000011001001111010", -- 12921 FREE #<CONS 0 12922>
 "00000000000000000011001001111011", -- 12922 FREE #<CONS 0 12923>
 "00000000000000000011001001111100", -- 12923 FREE #<CONS 0 12924>
 "00000000000000000011001001111101", -- 12924 FREE #<CONS 0 12925>
 "00000000000000000011001001111110", -- 12925 FREE #<CONS 0 12926>
 "00000000000000000011001001111111", -- 12926 FREE #<CONS 0 12927>
 "00000000000000000011001010000000", -- 12927 FREE #<CONS 0 12928>
 "00000000000000000011001010000001", -- 12928 FREE #<CONS 0 12929>
 "00000000000000000011001010000010", -- 12929 FREE #<CONS 0 12930>
 "00000000000000000011001010000011", -- 12930 FREE #<CONS 0 12931>
 "00000000000000000011001010000100", -- 12931 FREE #<CONS 0 12932>
 "00000000000000000011001010000101", -- 12932 FREE #<CONS 0 12933>
 "00000000000000000011001010000110", -- 12933 FREE #<CONS 0 12934>
 "00000000000000000011001010000111", -- 12934 FREE #<CONS 0 12935>
 "00000000000000000011001010001000", -- 12935 FREE #<CONS 0 12936>
 "00000000000000000011001010001001", -- 12936 FREE #<CONS 0 12937>
 "00000000000000000011001010001010", -- 12937 FREE #<CONS 0 12938>
 "00000000000000000011001010001011", -- 12938 FREE #<CONS 0 12939>
 "00000000000000000011001010001100", -- 12939 FREE #<CONS 0 12940>
 "00000000000000000011001010001101", -- 12940 FREE #<CONS 0 12941>
 "00000000000000000011001010001110", -- 12941 FREE #<CONS 0 12942>
 "00000000000000000011001010001111", -- 12942 FREE #<CONS 0 12943>
 "00000000000000000011001010010000", -- 12943 FREE #<CONS 0 12944>
 "00000000000000000011001010010001", -- 12944 FREE #<CONS 0 12945>
 "00000000000000000011001010010010", -- 12945 FREE #<CONS 0 12946>
 "00000000000000000011001010010011", -- 12946 FREE #<CONS 0 12947>
 "00000000000000000011001010010100", -- 12947 FREE #<CONS 0 12948>
 "00000000000000000011001010010101", -- 12948 FREE #<CONS 0 12949>
 "00000000000000000011001010010110", -- 12949 FREE #<CONS 0 12950>
 "00000000000000000011001010010111", -- 12950 FREE #<CONS 0 12951>
 "00000000000000000011001010011000", -- 12951 FREE #<CONS 0 12952>
 "00000000000000000011001010011001", -- 12952 FREE #<CONS 0 12953>
 "00000000000000000011001010011010", -- 12953 FREE #<CONS 0 12954>
 "00000000000000000011001010011011", -- 12954 FREE #<CONS 0 12955>
 "00000000000000000011001010011100", -- 12955 FREE #<CONS 0 12956>
 "00000000000000000011001010011101", -- 12956 FREE #<CONS 0 12957>
 "00000000000000000011001010011110", -- 12957 FREE #<CONS 0 12958>
 "00000000000000000011001010011111", -- 12958 FREE #<CONS 0 12959>
 "00000000000000000011001010100000", -- 12959 FREE #<CONS 0 12960>
 "00000000000000000011001010100001", -- 12960 FREE #<CONS 0 12961>
 "00000000000000000011001010100010", -- 12961 FREE #<CONS 0 12962>
 "00000000000000000011001010100011", -- 12962 FREE #<CONS 0 12963>
 "00000000000000000011001010100100", -- 12963 FREE #<CONS 0 12964>
 "00000000000000000011001010100101", -- 12964 FREE #<CONS 0 12965>
 "00000000000000000011001010100110", -- 12965 FREE #<CONS 0 12966>
 "00000000000000000011001010100111", -- 12966 FREE #<CONS 0 12967>
 "00000000000000000011001010101000", -- 12967 FREE #<CONS 0 12968>
 "00000000000000000011001010101001", -- 12968 FREE #<CONS 0 12969>
 "00000000000000000011001010101010", -- 12969 FREE #<CONS 0 12970>
 "00000000000000000011001010101011", -- 12970 FREE #<CONS 0 12971>
 "00000000000000000011001010101100", -- 12971 FREE #<CONS 0 12972>
 "00000000000000000011001010101101", -- 12972 FREE #<CONS 0 12973>
 "00000000000000000011001010101110", -- 12973 FREE #<CONS 0 12974>
 "00000000000000000011001010101111", -- 12974 FREE #<CONS 0 12975>
 "00000000000000000011001010110000", -- 12975 FREE #<CONS 0 12976>
 "00000000000000000011001010110001", -- 12976 FREE #<CONS 0 12977>
 "00000000000000000011001010110010", -- 12977 FREE #<CONS 0 12978>
 "00000000000000000011001010110011", -- 12978 FREE #<CONS 0 12979>
 "00000000000000000011001010110100", -- 12979 FREE #<CONS 0 12980>
 "00000000000000000011001010110101", -- 12980 FREE #<CONS 0 12981>
 "00000000000000000011001010110110", -- 12981 FREE #<CONS 0 12982>
 "00000000000000000011001010110111", -- 12982 FREE #<CONS 0 12983>
 "00000000000000000011001010111000", -- 12983 FREE #<CONS 0 12984>
 "00000000000000000011001010111001", -- 12984 FREE #<CONS 0 12985>
 "00000000000000000011001010111010", -- 12985 FREE #<CONS 0 12986>
 "00000000000000000011001010111011", -- 12986 FREE #<CONS 0 12987>
 "00000000000000000011001010111100", -- 12987 FREE #<CONS 0 12988>
 "00000000000000000011001010111101", -- 12988 FREE #<CONS 0 12989>
 "00000000000000000011001010111110", -- 12989 FREE #<CONS 0 12990>
 "00000000000000000011001010111111", -- 12990 FREE #<CONS 0 12991>
 "00000000000000000011001011000000", -- 12991 FREE #<CONS 0 12992>
 "00000000000000000011001011000001", -- 12992 FREE #<CONS 0 12993>
 "00000000000000000011001011000010", -- 12993 FREE #<CONS 0 12994>
 "00000000000000000011001011000011", -- 12994 FREE #<CONS 0 12995>
 "00000000000000000011001011000100", -- 12995 FREE #<CONS 0 12996>
 "00000000000000000011001011000101", -- 12996 FREE #<CONS 0 12997>
 "00000000000000000011001011000110", -- 12997 FREE #<CONS 0 12998>
 "00000000000000000011001011000111", -- 12998 FREE #<CONS 0 12999>
 "00000000000000000011001011001000", -- 12999 FREE #<CONS 0 13000>
 "00000000000000000011001011001001", -- 13000 FREE #<CONS 0 13001>
 "00000000000000000011001011001010", -- 13001 FREE #<CONS 0 13002>
 "00000000000000000011001011001011", -- 13002 FREE #<CONS 0 13003>
 "00000000000000000011001011001100", -- 13003 FREE #<CONS 0 13004>
 "00000000000000000011001011001101", -- 13004 FREE #<CONS 0 13005>
 "00000000000000000011001011001110", -- 13005 FREE #<CONS 0 13006>
 "00000000000000000011001011001111", -- 13006 FREE #<CONS 0 13007>
 "00000000000000000011001011010000", -- 13007 FREE #<CONS 0 13008>
 "00000000000000000011001011010001", -- 13008 FREE #<CONS 0 13009>
 "00000000000000000011001011010010", -- 13009 FREE #<CONS 0 13010>
 "00000000000000000011001011010011", -- 13010 FREE #<CONS 0 13011>
 "00000000000000000011001011010100", -- 13011 FREE #<CONS 0 13012>
 "00000000000000000011001011010101", -- 13012 FREE #<CONS 0 13013>
 "00000000000000000011001011010110", -- 13013 FREE #<CONS 0 13014>
 "00000000000000000011001011010111", -- 13014 FREE #<CONS 0 13015>
 "00000000000000000011001011011000", -- 13015 FREE #<CONS 0 13016>
 "00000000000000000011001011011001", -- 13016 FREE #<CONS 0 13017>
 "00000000000000000011001011011010", -- 13017 FREE #<CONS 0 13018>
 "00000000000000000011001011011011", -- 13018 FREE #<CONS 0 13019>
 "00000000000000000011001011011100", -- 13019 FREE #<CONS 0 13020>
 "00000000000000000011001011011101", -- 13020 FREE #<CONS 0 13021>
 "00000000000000000011001011011110", -- 13021 FREE #<CONS 0 13022>
 "00000000000000000011001011011111", -- 13022 FREE #<CONS 0 13023>
 "00000000000000000011001011100000", -- 13023 FREE #<CONS 0 13024>
 "00000000000000000011001011100001", -- 13024 FREE #<CONS 0 13025>
 "00000000000000000011001011100010", -- 13025 FREE #<CONS 0 13026>
 "00000000000000000011001011100011", -- 13026 FREE #<CONS 0 13027>
 "00000000000000000011001011100100", -- 13027 FREE #<CONS 0 13028>
 "00000000000000000011001011100101", -- 13028 FREE #<CONS 0 13029>
 "00000000000000000011001011100110", -- 13029 FREE #<CONS 0 13030>
 "00000000000000000011001011100111", -- 13030 FREE #<CONS 0 13031>
 "00000000000000000011001011101000", -- 13031 FREE #<CONS 0 13032>
 "00000000000000000011001011101001", -- 13032 FREE #<CONS 0 13033>
 "00000000000000000011001011101010", -- 13033 FREE #<CONS 0 13034>
 "00000000000000000011001011101011", -- 13034 FREE #<CONS 0 13035>
 "00000000000000000011001011101100", -- 13035 FREE #<CONS 0 13036>
 "00000000000000000011001011101101", -- 13036 FREE #<CONS 0 13037>
 "00000000000000000011001011101110", -- 13037 FREE #<CONS 0 13038>
 "00000000000000000011001011101111", -- 13038 FREE #<CONS 0 13039>
 "00000000000000000011001011110000", -- 13039 FREE #<CONS 0 13040>
 "00000000000000000011001011110001", -- 13040 FREE #<CONS 0 13041>
 "00000000000000000011001011110010", -- 13041 FREE #<CONS 0 13042>
 "00000000000000000011001011110011", -- 13042 FREE #<CONS 0 13043>
 "00000000000000000011001011110100", -- 13043 FREE #<CONS 0 13044>
 "00000000000000000011001011110101", -- 13044 FREE #<CONS 0 13045>
 "00000000000000000011001011110110", -- 13045 FREE #<CONS 0 13046>
 "00000000000000000011001011110111", -- 13046 FREE #<CONS 0 13047>
 "00000000000000000011001011111000", -- 13047 FREE #<CONS 0 13048>
 "00000000000000000011001011111001", -- 13048 FREE #<CONS 0 13049>
 "00000000000000000011001011111010", -- 13049 FREE #<CONS 0 13050>
 "00000000000000000011001011111011", -- 13050 FREE #<CONS 0 13051>
 "00000000000000000011001011111100", -- 13051 FREE #<CONS 0 13052>
 "00000000000000000011001011111101", -- 13052 FREE #<CONS 0 13053>
 "00000000000000000011001011111110", -- 13053 FREE #<CONS 0 13054>
 "00000000000000000011001011111111", -- 13054 FREE #<CONS 0 13055>
 "00000000000000000011001100000000", -- 13055 FREE #<CONS 0 13056>
 "00000000000000000011001100000001", -- 13056 FREE #<CONS 0 13057>
 "00000000000000000011001100000010", -- 13057 FREE #<CONS 0 13058>
 "00000000000000000011001100000011", -- 13058 FREE #<CONS 0 13059>
 "00000000000000000011001100000100", -- 13059 FREE #<CONS 0 13060>
 "00000000000000000011001100000101", -- 13060 FREE #<CONS 0 13061>
 "00000000000000000011001100000110", -- 13061 FREE #<CONS 0 13062>
 "00000000000000000011001100000111", -- 13062 FREE #<CONS 0 13063>
 "00000000000000000011001100001000", -- 13063 FREE #<CONS 0 13064>
 "00000000000000000011001100001001", -- 13064 FREE #<CONS 0 13065>
 "00000000000000000011001100001010", -- 13065 FREE #<CONS 0 13066>
 "00000000000000000011001100001011", -- 13066 FREE #<CONS 0 13067>
 "00000000000000000011001100001100", -- 13067 FREE #<CONS 0 13068>
 "00000000000000000011001100001101", -- 13068 FREE #<CONS 0 13069>
 "00000000000000000011001100001110", -- 13069 FREE #<CONS 0 13070>
 "00000000000000000011001100001111", -- 13070 FREE #<CONS 0 13071>
 "00000000000000000011001100010000", -- 13071 FREE #<CONS 0 13072>
 "00000000000000000011001100010001", -- 13072 FREE #<CONS 0 13073>
 "00000000000000000011001100010010", -- 13073 FREE #<CONS 0 13074>
 "00000000000000000011001100010011", -- 13074 FREE #<CONS 0 13075>
 "00000000000000000011001100010100", -- 13075 FREE #<CONS 0 13076>
 "00000000000000000011001100010101", -- 13076 FREE #<CONS 0 13077>
 "00000000000000000011001100010110", -- 13077 FREE #<CONS 0 13078>
 "00000000000000000011001100010111", -- 13078 FREE #<CONS 0 13079>
 "00000000000000000011001100011000", -- 13079 FREE #<CONS 0 13080>
 "00000000000000000011001100011001", -- 13080 FREE #<CONS 0 13081>
 "00000000000000000011001100011010", -- 13081 FREE #<CONS 0 13082>
 "00000000000000000011001100011011", -- 13082 FREE #<CONS 0 13083>
 "00000000000000000011001100011100", -- 13083 FREE #<CONS 0 13084>
 "00000000000000000011001100011101", -- 13084 FREE #<CONS 0 13085>
 "00000000000000000011001100011110", -- 13085 FREE #<CONS 0 13086>
 "00000000000000000011001100011111", -- 13086 FREE #<CONS 0 13087>
 "00000000000000000011001100100000", -- 13087 FREE #<CONS 0 13088>
 "00000000000000000011001100100001", -- 13088 FREE #<CONS 0 13089>
 "00000000000000000011001100100010", -- 13089 FREE #<CONS 0 13090>
 "00000000000000000011001100100011", -- 13090 FREE #<CONS 0 13091>
 "00000000000000000011001100100100", -- 13091 FREE #<CONS 0 13092>
 "00000000000000000011001100100101", -- 13092 FREE #<CONS 0 13093>
 "00000000000000000011001100100110", -- 13093 FREE #<CONS 0 13094>
 "00000000000000000011001100100111", -- 13094 FREE #<CONS 0 13095>
 "00000000000000000011001100101000", -- 13095 FREE #<CONS 0 13096>
 "00000000000000000011001100101001", -- 13096 FREE #<CONS 0 13097>
 "00000000000000000011001100101010", -- 13097 FREE #<CONS 0 13098>
 "00000000000000000011001100101011", -- 13098 FREE #<CONS 0 13099>
 "00000000000000000011001100101100", -- 13099 FREE #<CONS 0 13100>
 "00000000000000000011001100101101", -- 13100 FREE #<CONS 0 13101>
 "00000000000000000011001100101110", -- 13101 FREE #<CONS 0 13102>
 "00000000000000000011001100101111", -- 13102 FREE #<CONS 0 13103>
 "00000000000000000011001100110000", -- 13103 FREE #<CONS 0 13104>
 "00000000000000000011001100110001", -- 13104 FREE #<CONS 0 13105>
 "00000000000000000011001100110010", -- 13105 FREE #<CONS 0 13106>
 "00000000000000000011001100110011", -- 13106 FREE #<CONS 0 13107>
 "00000000000000000011001100110100", -- 13107 FREE #<CONS 0 13108>
 "00000000000000000011001100110101", -- 13108 FREE #<CONS 0 13109>
 "00000000000000000011001100110110", -- 13109 FREE #<CONS 0 13110>
 "00000000000000000011001100110111", -- 13110 FREE #<CONS 0 13111>
 "00000000000000000011001100111000", -- 13111 FREE #<CONS 0 13112>
 "00000000000000000011001100111001", -- 13112 FREE #<CONS 0 13113>
 "00000000000000000011001100111010", -- 13113 FREE #<CONS 0 13114>
 "00000000000000000011001100111011", -- 13114 FREE #<CONS 0 13115>
 "00000000000000000011001100111100", -- 13115 FREE #<CONS 0 13116>
 "00000000000000000011001100111101", -- 13116 FREE #<CONS 0 13117>
 "00000000000000000011001100111110", -- 13117 FREE #<CONS 0 13118>
 "00000000000000000011001100111111", -- 13118 FREE #<CONS 0 13119>
 "00000000000000000011001101000000", -- 13119 FREE #<CONS 0 13120>
 "00000000000000000011001101000001", -- 13120 FREE #<CONS 0 13121>
 "00000000000000000011001101000010", -- 13121 FREE #<CONS 0 13122>
 "00000000000000000011001101000011", -- 13122 FREE #<CONS 0 13123>
 "00000000000000000011001101000100", -- 13123 FREE #<CONS 0 13124>
 "00000000000000000011001101000101", -- 13124 FREE #<CONS 0 13125>
 "00000000000000000011001101000110", -- 13125 FREE #<CONS 0 13126>
 "00000000000000000011001101000111", -- 13126 FREE #<CONS 0 13127>
 "00000000000000000011001101001000", -- 13127 FREE #<CONS 0 13128>
 "00000000000000000011001101001001", -- 13128 FREE #<CONS 0 13129>
 "00000000000000000011001101001010", -- 13129 FREE #<CONS 0 13130>
 "00000000000000000011001101001011", -- 13130 FREE #<CONS 0 13131>
 "00000000000000000011001101001100", -- 13131 FREE #<CONS 0 13132>
 "00000000000000000011001101001101", -- 13132 FREE #<CONS 0 13133>
 "00000000000000000011001101001110", -- 13133 FREE #<CONS 0 13134>
 "00000000000000000011001101001111", -- 13134 FREE #<CONS 0 13135>
 "00000000000000000011001101010000", -- 13135 FREE #<CONS 0 13136>
 "00000000000000000011001101010001", -- 13136 FREE #<CONS 0 13137>
 "00000000000000000011001101010010", -- 13137 FREE #<CONS 0 13138>
 "00000000000000000011001101010011", -- 13138 FREE #<CONS 0 13139>
 "00000000000000000011001101010100", -- 13139 FREE #<CONS 0 13140>
 "00000000000000000011001101010101", -- 13140 FREE #<CONS 0 13141>
 "00000000000000000011001101010110", -- 13141 FREE #<CONS 0 13142>
 "00000000000000000011001101010111", -- 13142 FREE #<CONS 0 13143>
 "00000000000000000011001101011000", -- 13143 FREE #<CONS 0 13144>
 "00000000000000000011001101011001", -- 13144 FREE #<CONS 0 13145>
 "00000000000000000011001101011010", -- 13145 FREE #<CONS 0 13146>
 "00000000000000000011001101011011", -- 13146 FREE #<CONS 0 13147>
 "00000000000000000011001101011100", -- 13147 FREE #<CONS 0 13148>
 "00000000000000000011001101011101", -- 13148 FREE #<CONS 0 13149>
 "00000000000000000011001101011110", -- 13149 FREE #<CONS 0 13150>
 "00000000000000000011001101011111", -- 13150 FREE #<CONS 0 13151>
 "00000000000000000011001101100000", -- 13151 FREE #<CONS 0 13152>
 "00000000000000000011001101100001", -- 13152 FREE #<CONS 0 13153>
 "00000000000000000011001101100010", -- 13153 FREE #<CONS 0 13154>
 "00000000000000000011001101100011", -- 13154 FREE #<CONS 0 13155>
 "00000000000000000011001101100100", -- 13155 FREE #<CONS 0 13156>
 "00000000000000000011001101100101", -- 13156 FREE #<CONS 0 13157>
 "00000000000000000011001101100110", -- 13157 FREE #<CONS 0 13158>
 "00000000000000000011001101100111", -- 13158 FREE #<CONS 0 13159>
 "00000000000000000011001101101000", -- 13159 FREE #<CONS 0 13160>
 "00000000000000000011001101101001", -- 13160 FREE #<CONS 0 13161>
 "00000000000000000011001101101010", -- 13161 FREE #<CONS 0 13162>
 "00000000000000000011001101101011", -- 13162 FREE #<CONS 0 13163>
 "00000000000000000011001101101100", -- 13163 FREE #<CONS 0 13164>
 "00000000000000000011001101101101", -- 13164 FREE #<CONS 0 13165>
 "00000000000000000011001101101110", -- 13165 FREE #<CONS 0 13166>
 "00000000000000000011001101101111", -- 13166 FREE #<CONS 0 13167>
 "00000000000000000011001101110000", -- 13167 FREE #<CONS 0 13168>
 "00000000000000000011001101110001", -- 13168 FREE #<CONS 0 13169>
 "00000000000000000011001101110010", -- 13169 FREE #<CONS 0 13170>
 "00000000000000000011001101110011", -- 13170 FREE #<CONS 0 13171>
 "00000000000000000011001101110100", -- 13171 FREE #<CONS 0 13172>
 "00000000000000000011001101110101", -- 13172 FREE #<CONS 0 13173>
 "00000000000000000011001101110110", -- 13173 FREE #<CONS 0 13174>
 "00000000000000000011001101110111", -- 13174 FREE #<CONS 0 13175>
 "00000000000000000011001101111000", -- 13175 FREE #<CONS 0 13176>
 "00000000000000000011001101111001", -- 13176 FREE #<CONS 0 13177>
 "00000000000000000011001101111010", -- 13177 FREE #<CONS 0 13178>
 "00000000000000000011001101111011", -- 13178 FREE #<CONS 0 13179>
 "00000000000000000011001101111100", -- 13179 FREE #<CONS 0 13180>
 "00000000000000000011001101111101", -- 13180 FREE #<CONS 0 13181>
 "00000000000000000011001101111110", -- 13181 FREE #<CONS 0 13182>
 "00000000000000000011001101111111", -- 13182 FREE #<CONS 0 13183>
 "00000000000000000011001110000000", -- 13183 FREE #<CONS 0 13184>
 "00000000000000000011001110000001", -- 13184 FREE #<CONS 0 13185>
 "00000000000000000011001110000010", -- 13185 FREE #<CONS 0 13186>
 "00000000000000000011001110000011", -- 13186 FREE #<CONS 0 13187>
 "00000000000000000011001110000100", -- 13187 FREE #<CONS 0 13188>
 "00000000000000000011001110000101", -- 13188 FREE #<CONS 0 13189>
 "00000000000000000011001110000110", -- 13189 FREE #<CONS 0 13190>
 "00000000000000000011001110000111", -- 13190 FREE #<CONS 0 13191>
 "00000000000000000011001110001000", -- 13191 FREE #<CONS 0 13192>
 "00000000000000000011001110001001", -- 13192 FREE #<CONS 0 13193>
 "00000000000000000011001110001010", -- 13193 FREE #<CONS 0 13194>
 "00000000000000000011001110001011", -- 13194 FREE #<CONS 0 13195>
 "00000000000000000011001110001100", -- 13195 FREE #<CONS 0 13196>
 "00000000000000000011001110001101", -- 13196 FREE #<CONS 0 13197>
 "00000000000000000011001110001110", -- 13197 FREE #<CONS 0 13198>
 "00000000000000000011001110001111", -- 13198 FREE #<CONS 0 13199>
 "00000000000000000011001110010000", -- 13199 FREE #<CONS 0 13200>
 "00000000000000000011001110010001", -- 13200 FREE #<CONS 0 13201>
 "00000000000000000011001110010010", -- 13201 FREE #<CONS 0 13202>
 "00000000000000000011001110010011", -- 13202 FREE #<CONS 0 13203>
 "00000000000000000011001110010100", -- 13203 FREE #<CONS 0 13204>
 "00000000000000000011001110010101", -- 13204 FREE #<CONS 0 13205>
 "00000000000000000011001110010110", -- 13205 FREE #<CONS 0 13206>
 "00000000000000000011001110010111", -- 13206 FREE #<CONS 0 13207>
 "00000000000000000011001110011000", -- 13207 FREE #<CONS 0 13208>
 "00000000000000000011001110011001", -- 13208 FREE #<CONS 0 13209>
 "00000000000000000011001110011010", -- 13209 FREE #<CONS 0 13210>
 "00000000000000000011001110011011", -- 13210 FREE #<CONS 0 13211>
 "00000000000000000011001110011100", -- 13211 FREE #<CONS 0 13212>
 "00000000000000000011001110011101", -- 13212 FREE #<CONS 0 13213>
 "00000000000000000011001110011110", -- 13213 FREE #<CONS 0 13214>
 "00000000000000000011001110011111", -- 13214 FREE #<CONS 0 13215>
 "00000000000000000011001110100000", -- 13215 FREE #<CONS 0 13216>
 "00000000000000000011001110100001", -- 13216 FREE #<CONS 0 13217>
 "00000000000000000011001110100010", -- 13217 FREE #<CONS 0 13218>
 "00000000000000000011001110100011", -- 13218 FREE #<CONS 0 13219>
 "00000000000000000011001110100100", -- 13219 FREE #<CONS 0 13220>
 "00000000000000000011001110100101", -- 13220 FREE #<CONS 0 13221>
 "00000000000000000011001110100110", -- 13221 FREE #<CONS 0 13222>
 "00000000000000000011001110100111", -- 13222 FREE #<CONS 0 13223>
 "00000000000000000011001110101000", -- 13223 FREE #<CONS 0 13224>
 "00000000000000000011001110101001", -- 13224 FREE #<CONS 0 13225>
 "00000000000000000011001110101010", -- 13225 FREE #<CONS 0 13226>
 "00000000000000000011001110101011", -- 13226 FREE #<CONS 0 13227>
 "00000000000000000011001110101100", -- 13227 FREE #<CONS 0 13228>
 "00000000000000000011001110101101", -- 13228 FREE #<CONS 0 13229>
 "00000000000000000011001110101110", -- 13229 FREE #<CONS 0 13230>
 "00000000000000000011001110101111", -- 13230 FREE #<CONS 0 13231>
 "00000000000000000011001110110000", -- 13231 FREE #<CONS 0 13232>
 "00000000000000000011001110110001", -- 13232 FREE #<CONS 0 13233>
 "00000000000000000011001110110010", -- 13233 FREE #<CONS 0 13234>
 "00000000000000000011001110110011", -- 13234 FREE #<CONS 0 13235>
 "00000000000000000011001110110100", -- 13235 FREE #<CONS 0 13236>
 "00000000000000000011001110110101", -- 13236 FREE #<CONS 0 13237>
 "00000000000000000011001110110110", -- 13237 FREE #<CONS 0 13238>
 "00000000000000000011001110110111", -- 13238 FREE #<CONS 0 13239>
 "00000000000000000011001110111000", -- 13239 FREE #<CONS 0 13240>
 "00000000000000000011001110111001", -- 13240 FREE #<CONS 0 13241>
 "00000000000000000011001110111010", -- 13241 FREE #<CONS 0 13242>
 "00000000000000000011001110111011", -- 13242 FREE #<CONS 0 13243>
 "00000000000000000011001110111100", -- 13243 FREE #<CONS 0 13244>
 "00000000000000000011001110111101", -- 13244 FREE #<CONS 0 13245>
 "00000000000000000011001110111110", -- 13245 FREE #<CONS 0 13246>
 "00000000000000000011001110111111", -- 13246 FREE #<CONS 0 13247>
 "00000000000000000011001111000000", -- 13247 FREE #<CONS 0 13248>
 "00000000000000000011001111000001", -- 13248 FREE #<CONS 0 13249>
 "00000000000000000011001111000010", -- 13249 FREE #<CONS 0 13250>
 "00000000000000000011001111000011", -- 13250 FREE #<CONS 0 13251>
 "00000000000000000011001111000100", -- 13251 FREE #<CONS 0 13252>
 "00000000000000000011001111000101", -- 13252 FREE #<CONS 0 13253>
 "00000000000000000011001111000110", -- 13253 FREE #<CONS 0 13254>
 "00000000000000000011001111000111", -- 13254 FREE #<CONS 0 13255>
 "00000000000000000011001111001000", -- 13255 FREE #<CONS 0 13256>
 "00000000000000000011001111001001", -- 13256 FREE #<CONS 0 13257>
 "00000000000000000011001111001010", -- 13257 FREE #<CONS 0 13258>
 "00000000000000000011001111001011", -- 13258 FREE #<CONS 0 13259>
 "00000000000000000011001111001100", -- 13259 FREE #<CONS 0 13260>
 "00000000000000000011001111001101", -- 13260 FREE #<CONS 0 13261>
 "00000000000000000011001111001110", -- 13261 FREE #<CONS 0 13262>
 "00000000000000000011001111001111", -- 13262 FREE #<CONS 0 13263>
 "00000000000000000011001111010000", -- 13263 FREE #<CONS 0 13264>
 "00000000000000000011001111010001", -- 13264 FREE #<CONS 0 13265>
 "00000000000000000011001111010010", -- 13265 FREE #<CONS 0 13266>
 "00000000000000000011001111010011", -- 13266 FREE #<CONS 0 13267>
 "00000000000000000011001111010100", -- 13267 FREE #<CONS 0 13268>
 "00000000000000000011001111010101", -- 13268 FREE #<CONS 0 13269>
 "00000000000000000011001111010110", -- 13269 FREE #<CONS 0 13270>
 "00000000000000000011001111010111", -- 13270 FREE #<CONS 0 13271>
 "00000000000000000011001111011000", -- 13271 FREE #<CONS 0 13272>
 "00000000000000000011001111011001", -- 13272 FREE #<CONS 0 13273>
 "00000000000000000011001111011010", -- 13273 FREE #<CONS 0 13274>
 "00000000000000000011001111011011", -- 13274 FREE #<CONS 0 13275>
 "00000000000000000011001111011100", -- 13275 FREE #<CONS 0 13276>
 "00000000000000000011001111011101", -- 13276 FREE #<CONS 0 13277>
 "00000000000000000011001111011110", -- 13277 FREE #<CONS 0 13278>
 "00000000000000000011001111011111", -- 13278 FREE #<CONS 0 13279>
 "00000000000000000011001111100000", -- 13279 FREE #<CONS 0 13280>
 "00000000000000000011001111100001", -- 13280 FREE #<CONS 0 13281>
 "00000000000000000011001111100010", -- 13281 FREE #<CONS 0 13282>
 "00000000000000000011001111100011", -- 13282 FREE #<CONS 0 13283>
 "00000000000000000011001111100100", -- 13283 FREE #<CONS 0 13284>
 "00000000000000000011001111100101", -- 13284 FREE #<CONS 0 13285>
 "00000000000000000011001111100110", -- 13285 FREE #<CONS 0 13286>
 "00000000000000000011001111100111", -- 13286 FREE #<CONS 0 13287>
 "00000000000000000011001111101000", -- 13287 FREE #<CONS 0 13288>
 "00000000000000000011001111101001", -- 13288 FREE #<CONS 0 13289>
 "00000000000000000011001111101010", -- 13289 FREE #<CONS 0 13290>
 "00000000000000000011001111101011", -- 13290 FREE #<CONS 0 13291>
 "00000000000000000011001111101100", -- 13291 FREE #<CONS 0 13292>
 "00000000000000000011001111101101", -- 13292 FREE #<CONS 0 13293>
 "00000000000000000011001111101110", -- 13293 FREE #<CONS 0 13294>
 "00000000000000000011001111101111", -- 13294 FREE #<CONS 0 13295>
 "00000000000000000011001111110000", -- 13295 FREE #<CONS 0 13296>
 "00000000000000000011001111110001", -- 13296 FREE #<CONS 0 13297>
 "00000000000000000011001111110010", -- 13297 FREE #<CONS 0 13298>
 "00000000000000000011001111110011", -- 13298 FREE #<CONS 0 13299>
 "00000000000000000011001111110100", -- 13299 FREE #<CONS 0 13300>
 "00000000000000000011001111110101", -- 13300 FREE #<CONS 0 13301>
 "00000000000000000011001111110110", -- 13301 FREE #<CONS 0 13302>
 "00000000000000000011001111110111", -- 13302 FREE #<CONS 0 13303>
 "00000000000000000011001111111000", -- 13303 FREE #<CONS 0 13304>
 "00000000000000000011001111111001", -- 13304 FREE #<CONS 0 13305>
 "00000000000000000011001111111010", -- 13305 FREE #<CONS 0 13306>
 "00000000000000000011001111111011", -- 13306 FREE #<CONS 0 13307>
 "00000000000000000011001111111100", -- 13307 FREE #<CONS 0 13308>
 "00000000000000000011001111111101", -- 13308 FREE #<CONS 0 13309>
 "00000000000000000011001111111110", -- 13309 FREE #<CONS 0 13310>
 "00000000000000000011001111111111", -- 13310 FREE #<CONS 0 13311>
 "00000000000000000011010000000000", -- 13311 FREE #<CONS 0 13312>
 "00000000000000000011010000000001", -- 13312 FREE #<CONS 0 13313>
 "00000000000000000011010000000010", -- 13313 FREE #<CONS 0 13314>
 "00000000000000000011010000000011", -- 13314 FREE #<CONS 0 13315>
 "00000000000000000011010000000100", -- 13315 FREE #<CONS 0 13316>
 "00000000000000000011010000000101", -- 13316 FREE #<CONS 0 13317>
 "00000000000000000011010000000110", -- 13317 FREE #<CONS 0 13318>
 "00000000000000000011010000000111", -- 13318 FREE #<CONS 0 13319>
 "00000000000000000011010000001000", -- 13319 FREE #<CONS 0 13320>
 "00000000000000000011010000001001", -- 13320 FREE #<CONS 0 13321>
 "00000000000000000011010000001010", -- 13321 FREE #<CONS 0 13322>
 "00000000000000000011010000001011", -- 13322 FREE #<CONS 0 13323>
 "00000000000000000011010000001100", -- 13323 FREE #<CONS 0 13324>
 "00000000000000000011010000001101", -- 13324 FREE #<CONS 0 13325>
 "00000000000000000011010000001110", -- 13325 FREE #<CONS 0 13326>
 "00000000000000000011010000001111", -- 13326 FREE #<CONS 0 13327>
 "00000000000000000011010000010000", -- 13327 FREE #<CONS 0 13328>
 "00000000000000000011010000010001", -- 13328 FREE #<CONS 0 13329>
 "00000000000000000011010000010010", -- 13329 FREE #<CONS 0 13330>
 "00000000000000000011010000010011", -- 13330 FREE #<CONS 0 13331>
 "00000000000000000011010000010100", -- 13331 FREE #<CONS 0 13332>
 "00000000000000000011010000010101", -- 13332 FREE #<CONS 0 13333>
 "00000000000000000011010000010110", -- 13333 FREE #<CONS 0 13334>
 "00000000000000000011010000010111", -- 13334 FREE #<CONS 0 13335>
 "00000000000000000011010000011000", -- 13335 FREE #<CONS 0 13336>
 "00000000000000000011010000011001", -- 13336 FREE #<CONS 0 13337>
 "00000000000000000011010000011010", -- 13337 FREE #<CONS 0 13338>
 "00000000000000000011010000011011", -- 13338 FREE #<CONS 0 13339>
 "00000000000000000011010000011100", -- 13339 FREE #<CONS 0 13340>
 "00000000000000000011010000011101", -- 13340 FREE #<CONS 0 13341>
 "00000000000000000011010000011110", -- 13341 FREE #<CONS 0 13342>
 "00000000000000000011010000011111", -- 13342 FREE #<CONS 0 13343>
 "00000000000000000011010000100000", -- 13343 FREE #<CONS 0 13344>
 "00000000000000000011010000100001", -- 13344 FREE #<CONS 0 13345>
 "00000000000000000011010000100010", -- 13345 FREE #<CONS 0 13346>
 "00000000000000000011010000100011", -- 13346 FREE #<CONS 0 13347>
 "00000000000000000011010000100100", -- 13347 FREE #<CONS 0 13348>
 "00000000000000000011010000100101", -- 13348 FREE #<CONS 0 13349>
 "00000000000000000011010000100110", -- 13349 FREE #<CONS 0 13350>
 "00000000000000000011010000100111", -- 13350 FREE #<CONS 0 13351>
 "00000000000000000011010000101000", -- 13351 FREE #<CONS 0 13352>
 "00000000000000000011010000101001", -- 13352 FREE #<CONS 0 13353>
 "00000000000000000011010000101010", -- 13353 FREE #<CONS 0 13354>
 "00000000000000000011010000101011", -- 13354 FREE #<CONS 0 13355>
 "00000000000000000011010000101100", -- 13355 FREE #<CONS 0 13356>
 "00000000000000000011010000101101", -- 13356 FREE #<CONS 0 13357>
 "00000000000000000011010000101110", -- 13357 FREE #<CONS 0 13358>
 "00000000000000000011010000101111", -- 13358 FREE #<CONS 0 13359>
 "00000000000000000011010000110000", -- 13359 FREE #<CONS 0 13360>
 "00000000000000000011010000110001", -- 13360 FREE #<CONS 0 13361>
 "00000000000000000011010000110010", -- 13361 FREE #<CONS 0 13362>
 "00000000000000000011010000110011", -- 13362 FREE #<CONS 0 13363>
 "00000000000000000011010000110100", -- 13363 FREE #<CONS 0 13364>
 "00000000000000000011010000110101", -- 13364 FREE #<CONS 0 13365>
 "00000000000000000011010000110110", -- 13365 FREE #<CONS 0 13366>
 "00000000000000000011010000110111", -- 13366 FREE #<CONS 0 13367>
 "00000000000000000011010000111000", -- 13367 FREE #<CONS 0 13368>
 "00000000000000000011010000111001", -- 13368 FREE #<CONS 0 13369>
 "00000000000000000011010000111010", -- 13369 FREE #<CONS 0 13370>
 "00000000000000000011010000111011", -- 13370 FREE #<CONS 0 13371>
 "00000000000000000011010000111100", -- 13371 FREE #<CONS 0 13372>
 "00000000000000000011010000111101", -- 13372 FREE #<CONS 0 13373>
 "00000000000000000011010000111110", -- 13373 FREE #<CONS 0 13374>
 "00000000000000000011010000111111", -- 13374 FREE #<CONS 0 13375>
 "00000000000000000011010001000000", -- 13375 FREE #<CONS 0 13376>
 "00000000000000000011010001000001", -- 13376 FREE #<CONS 0 13377>
 "00000000000000000011010001000010", -- 13377 FREE #<CONS 0 13378>
 "00000000000000000011010001000011", -- 13378 FREE #<CONS 0 13379>
 "00000000000000000011010001000100", -- 13379 FREE #<CONS 0 13380>
 "00000000000000000011010001000101", -- 13380 FREE #<CONS 0 13381>
 "00000000000000000011010001000110", -- 13381 FREE #<CONS 0 13382>
 "00000000000000000011010001000111", -- 13382 FREE #<CONS 0 13383>
 "00000000000000000011010001001000", -- 13383 FREE #<CONS 0 13384>
 "00000000000000000011010001001001", -- 13384 FREE #<CONS 0 13385>
 "00000000000000000011010001001010", -- 13385 FREE #<CONS 0 13386>
 "00000000000000000011010001001011", -- 13386 FREE #<CONS 0 13387>
 "00000000000000000011010001001100", -- 13387 FREE #<CONS 0 13388>
 "00000000000000000011010001001101", -- 13388 FREE #<CONS 0 13389>
 "00000000000000000011010001001110", -- 13389 FREE #<CONS 0 13390>
 "00000000000000000011010001001111", -- 13390 FREE #<CONS 0 13391>
 "00000000000000000011010001010000", -- 13391 FREE #<CONS 0 13392>
 "00000000000000000011010001010001", -- 13392 FREE #<CONS 0 13393>
 "00000000000000000011010001010010", -- 13393 FREE #<CONS 0 13394>
 "00000000000000000011010001010011", -- 13394 FREE #<CONS 0 13395>
 "00000000000000000011010001010100", -- 13395 FREE #<CONS 0 13396>
 "00000000000000000011010001010101", -- 13396 FREE #<CONS 0 13397>
 "00000000000000000011010001010110", -- 13397 FREE #<CONS 0 13398>
 "00000000000000000011010001010111", -- 13398 FREE #<CONS 0 13399>
 "00000000000000000011010001011000", -- 13399 FREE #<CONS 0 13400>
 "00000000000000000011010001011001", -- 13400 FREE #<CONS 0 13401>
 "00000000000000000011010001011010", -- 13401 FREE #<CONS 0 13402>
 "00000000000000000011010001011011", -- 13402 FREE #<CONS 0 13403>
 "00000000000000000011010001011100", -- 13403 FREE #<CONS 0 13404>
 "00000000000000000011010001011101", -- 13404 FREE #<CONS 0 13405>
 "00000000000000000011010001011110", -- 13405 FREE #<CONS 0 13406>
 "00000000000000000011010001011111", -- 13406 FREE #<CONS 0 13407>
 "00000000000000000011010001100000", -- 13407 FREE #<CONS 0 13408>
 "00000000000000000011010001100001", -- 13408 FREE #<CONS 0 13409>
 "00000000000000000011010001100010", -- 13409 FREE #<CONS 0 13410>
 "00000000000000000011010001100011", -- 13410 FREE #<CONS 0 13411>
 "00000000000000000011010001100100", -- 13411 FREE #<CONS 0 13412>
 "00000000000000000011010001100101", -- 13412 FREE #<CONS 0 13413>
 "00000000000000000011010001100110", -- 13413 FREE #<CONS 0 13414>
 "00000000000000000011010001100111", -- 13414 FREE #<CONS 0 13415>
 "00000000000000000011010001101000", -- 13415 FREE #<CONS 0 13416>
 "00000000000000000011010001101001", -- 13416 FREE #<CONS 0 13417>
 "00000000000000000011010001101010", -- 13417 FREE #<CONS 0 13418>
 "00000000000000000011010001101011", -- 13418 FREE #<CONS 0 13419>
 "00000000000000000011010001101100", -- 13419 FREE #<CONS 0 13420>
 "00000000000000000011010001101101", -- 13420 FREE #<CONS 0 13421>
 "00000000000000000011010001101110", -- 13421 FREE #<CONS 0 13422>
 "00000000000000000011010001101111", -- 13422 FREE #<CONS 0 13423>
 "00000000000000000011010001110000", -- 13423 FREE #<CONS 0 13424>
 "00000000000000000011010001110001", -- 13424 FREE #<CONS 0 13425>
 "00000000000000000011010001110010", -- 13425 FREE #<CONS 0 13426>
 "00000000000000000011010001110011", -- 13426 FREE #<CONS 0 13427>
 "00000000000000000011010001110100", -- 13427 FREE #<CONS 0 13428>
 "00000000000000000011010001110101", -- 13428 FREE #<CONS 0 13429>
 "00000000000000000011010001110110", -- 13429 FREE #<CONS 0 13430>
 "00000000000000000011010001110111", -- 13430 FREE #<CONS 0 13431>
 "00000000000000000011010001111000", -- 13431 FREE #<CONS 0 13432>
 "00000000000000000011010001111001", -- 13432 FREE #<CONS 0 13433>
 "00000000000000000011010001111010", -- 13433 FREE #<CONS 0 13434>
 "00000000000000000011010001111011", -- 13434 FREE #<CONS 0 13435>
 "00000000000000000011010001111100", -- 13435 FREE #<CONS 0 13436>
 "00000000000000000011010001111101", -- 13436 FREE #<CONS 0 13437>
 "00000000000000000011010001111110", -- 13437 FREE #<CONS 0 13438>
 "00000000000000000011010001111111", -- 13438 FREE #<CONS 0 13439>
 "00000000000000000011010010000000", -- 13439 FREE #<CONS 0 13440>
 "00000000000000000011010010000001", -- 13440 FREE #<CONS 0 13441>
 "00000000000000000011010010000010", -- 13441 FREE #<CONS 0 13442>
 "00000000000000000011010010000011", -- 13442 FREE #<CONS 0 13443>
 "00000000000000000011010010000100", -- 13443 FREE #<CONS 0 13444>
 "00000000000000000011010010000101", -- 13444 FREE #<CONS 0 13445>
 "00000000000000000011010010000110", -- 13445 FREE #<CONS 0 13446>
 "00000000000000000011010010000111", -- 13446 FREE #<CONS 0 13447>
 "00000000000000000011010010001000", -- 13447 FREE #<CONS 0 13448>
 "00000000000000000011010010001001", -- 13448 FREE #<CONS 0 13449>
 "00000000000000000011010010001010", -- 13449 FREE #<CONS 0 13450>
 "00000000000000000011010010001011", -- 13450 FREE #<CONS 0 13451>
 "00000000000000000011010010001100", -- 13451 FREE #<CONS 0 13452>
 "00000000000000000011010010001101", -- 13452 FREE #<CONS 0 13453>
 "00000000000000000011010010001110", -- 13453 FREE #<CONS 0 13454>
 "00000000000000000011010010001111", -- 13454 FREE #<CONS 0 13455>
 "00000000000000000011010010010000", -- 13455 FREE #<CONS 0 13456>
 "00000000000000000011010010010001", -- 13456 FREE #<CONS 0 13457>
 "00000000000000000011010010010010", -- 13457 FREE #<CONS 0 13458>
 "00000000000000000011010010010011", -- 13458 FREE #<CONS 0 13459>
 "00000000000000000011010010010100", -- 13459 FREE #<CONS 0 13460>
 "00000000000000000011010010010101", -- 13460 FREE #<CONS 0 13461>
 "00000000000000000011010010010110", -- 13461 FREE #<CONS 0 13462>
 "00000000000000000011010010010111", -- 13462 FREE #<CONS 0 13463>
 "00000000000000000011010010011000", -- 13463 FREE #<CONS 0 13464>
 "00000000000000000011010010011001", -- 13464 FREE #<CONS 0 13465>
 "00000000000000000011010010011010", -- 13465 FREE #<CONS 0 13466>
 "00000000000000000011010010011011", -- 13466 FREE #<CONS 0 13467>
 "00000000000000000011010010011100", -- 13467 FREE #<CONS 0 13468>
 "00000000000000000011010010011101", -- 13468 FREE #<CONS 0 13469>
 "00000000000000000011010010011110", -- 13469 FREE #<CONS 0 13470>
 "00000000000000000011010010011111", -- 13470 FREE #<CONS 0 13471>
 "00000000000000000011010010100000", -- 13471 FREE #<CONS 0 13472>
 "00000000000000000011010010100001", -- 13472 FREE #<CONS 0 13473>
 "00000000000000000011010010100010", -- 13473 FREE #<CONS 0 13474>
 "00000000000000000011010010100011", -- 13474 FREE #<CONS 0 13475>
 "00000000000000000011010010100100", -- 13475 FREE #<CONS 0 13476>
 "00000000000000000011010010100101", -- 13476 FREE #<CONS 0 13477>
 "00000000000000000011010010100110", -- 13477 FREE #<CONS 0 13478>
 "00000000000000000011010010100111", -- 13478 FREE #<CONS 0 13479>
 "00000000000000000011010010101000", -- 13479 FREE #<CONS 0 13480>
 "00000000000000000011010010101001", -- 13480 FREE #<CONS 0 13481>
 "00000000000000000011010010101010", -- 13481 FREE #<CONS 0 13482>
 "00000000000000000011010010101011", -- 13482 FREE #<CONS 0 13483>
 "00000000000000000011010010101100", -- 13483 FREE #<CONS 0 13484>
 "00000000000000000011010010101101", -- 13484 FREE #<CONS 0 13485>
 "00000000000000000011010010101110", -- 13485 FREE #<CONS 0 13486>
 "00000000000000000011010010101111", -- 13486 FREE #<CONS 0 13487>
 "00000000000000000011010010110000", -- 13487 FREE #<CONS 0 13488>
 "00000000000000000011010010110001", -- 13488 FREE #<CONS 0 13489>
 "00000000000000000011010010110010", -- 13489 FREE #<CONS 0 13490>
 "00000000000000000011010010110011", -- 13490 FREE #<CONS 0 13491>
 "00000000000000000011010010110100", -- 13491 FREE #<CONS 0 13492>
 "00000000000000000011010010110101", -- 13492 FREE #<CONS 0 13493>
 "00000000000000000011010010110110", -- 13493 FREE #<CONS 0 13494>
 "00000000000000000011010010110111", -- 13494 FREE #<CONS 0 13495>
 "00000000000000000011010010111000", -- 13495 FREE #<CONS 0 13496>
 "00000000000000000011010010111001", -- 13496 FREE #<CONS 0 13497>
 "00000000000000000011010010111010", -- 13497 FREE #<CONS 0 13498>
 "00000000000000000011010010111011", -- 13498 FREE #<CONS 0 13499>
 "00000000000000000011010010111100", -- 13499 FREE #<CONS 0 13500>
 "00000000000000000011010010111101", -- 13500 FREE #<CONS 0 13501>
 "00000000000000000011010010111110", -- 13501 FREE #<CONS 0 13502>
 "00000000000000000011010010111111", -- 13502 FREE #<CONS 0 13503>
 "00000000000000000011010011000000", -- 13503 FREE #<CONS 0 13504>
 "00000000000000000011010011000001", -- 13504 FREE #<CONS 0 13505>
 "00000000000000000011010011000010", -- 13505 FREE #<CONS 0 13506>
 "00000000000000000011010011000011", -- 13506 FREE #<CONS 0 13507>
 "00000000000000000011010011000100", -- 13507 FREE #<CONS 0 13508>
 "00000000000000000011010011000101", -- 13508 FREE #<CONS 0 13509>
 "00000000000000000011010011000110", -- 13509 FREE #<CONS 0 13510>
 "00000000000000000011010011000111", -- 13510 FREE #<CONS 0 13511>
 "00000000000000000011010011001000", -- 13511 FREE #<CONS 0 13512>
 "00000000000000000011010011001001", -- 13512 FREE #<CONS 0 13513>
 "00000000000000000011010011001010", -- 13513 FREE #<CONS 0 13514>
 "00000000000000000011010011001011", -- 13514 FREE #<CONS 0 13515>
 "00000000000000000011010011001100", -- 13515 FREE #<CONS 0 13516>
 "00000000000000000011010011001101", -- 13516 FREE #<CONS 0 13517>
 "00000000000000000011010011001110", -- 13517 FREE #<CONS 0 13518>
 "00000000000000000011010011001111", -- 13518 FREE #<CONS 0 13519>
 "00000000000000000011010011010000", -- 13519 FREE #<CONS 0 13520>
 "00000000000000000011010011010001", -- 13520 FREE #<CONS 0 13521>
 "00000000000000000011010011010010", -- 13521 FREE #<CONS 0 13522>
 "00000000000000000011010011010011", -- 13522 FREE #<CONS 0 13523>
 "00000000000000000011010011010100", -- 13523 FREE #<CONS 0 13524>
 "00000000000000000011010011010101", -- 13524 FREE #<CONS 0 13525>
 "00000000000000000011010011010110", -- 13525 FREE #<CONS 0 13526>
 "00000000000000000011010011010111", -- 13526 FREE #<CONS 0 13527>
 "00000000000000000011010011011000", -- 13527 FREE #<CONS 0 13528>
 "00000000000000000011010011011001", -- 13528 FREE #<CONS 0 13529>
 "00000000000000000011010011011010", -- 13529 FREE #<CONS 0 13530>
 "00000000000000000011010011011011", -- 13530 FREE #<CONS 0 13531>
 "00000000000000000011010011011100", -- 13531 FREE #<CONS 0 13532>
 "00000000000000000011010011011101", -- 13532 FREE #<CONS 0 13533>
 "00000000000000000011010011011110", -- 13533 FREE #<CONS 0 13534>
 "00000000000000000011010011011111", -- 13534 FREE #<CONS 0 13535>
 "00000000000000000011010011100000", -- 13535 FREE #<CONS 0 13536>
 "00000000000000000011010011100001", -- 13536 FREE #<CONS 0 13537>
 "00000000000000000011010011100010", -- 13537 FREE #<CONS 0 13538>
 "00000000000000000011010011100011", -- 13538 FREE #<CONS 0 13539>
 "00000000000000000011010011100100", -- 13539 FREE #<CONS 0 13540>
 "00000000000000000011010011100101", -- 13540 FREE #<CONS 0 13541>
 "00000000000000000011010011100110", -- 13541 FREE #<CONS 0 13542>
 "00000000000000000011010011100111", -- 13542 FREE #<CONS 0 13543>
 "00000000000000000011010011101000", -- 13543 FREE #<CONS 0 13544>
 "00000000000000000011010011101001", -- 13544 FREE #<CONS 0 13545>
 "00000000000000000011010011101010", -- 13545 FREE #<CONS 0 13546>
 "00000000000000000011010011101011", -- 13546 FREE #<CONS 0 13547>
 "00000000000000000011010011101100", -- 13547 FREE #<CONS 0 13548>
 "00000000000000000011010011101101", -- 13548 FREE #<CONS 0 13549>
 "00000000000000000011010011101110", -- 13549 FREE #<CONS 0 13550>
 "00000000000000000011010011101111", -- 13550 FREE #<CONS 0 13551>
 "00000000000000000011010011110000", -- 13551 FREE #<CONS 0 13552>
 "00000000000000000011010011110001", -- 13552 FREE #<CONS 0 13553>
 "00000000000000000011010011110010", -- 13553 FREE #<CONS 0 13554>
 "00000000000000000011010011110011", -- 13554 FREE #<CONS 0 13555>
 "00000000000000000011010011110100", -- 13555 FREE #<CONS 0 13556>
 "00000000000000000011010011110101", -- 13556 FREE #<CONS 0 13557>
 "00000000000000000011010011110110", -- 13557 FREE #<CONS 0 13558>
 "00000000000000000011010011110111", -- 13558 FREE #<CONS 0 13559>
 "00000000000000000011010011111000", -- 13559 FREE #<CONS 0 13560>
 "00000000000000000011010011111001", -- 13560 FREE #<CONS 0 13561>
 "00000000000000000011010011111010", -- 13561 FREE #<CONS 0 13562>
 "00000000000000000011010011111011", -- 13562 FREE #<CONS 0 13563>
 "00000000000000000011010011111100", -- 13563 FREE #<CONS 0 13564>
 "00000000000000000011010011111101", -- 13564 FREE #<CONS 0 13565>
 "00000000000000000011010011111110", -- 13565 FREE #<CONS 0 13566>
 "00000000000000000011010011111111", -- 13566 FREE #<CONS 0 13567>
 "00000000000000000011010100000000", -- 13567 FREE #<CONS 0 13568>
 "00000000000000000011010100000001", -- 13568 FREE #<CONS 0 13569>
 "00000000000000000011010100000010", -- 13569 FREE #<CONS 0 13570>
 "00000000000000000011010100000011", -- 13570 FREE #<CONS 0 13571>
 "00000000000000000011010100000100", -- 13571 FREE #<CONS 0 13572>
 "00000000000000000011010100000101", -- 13572 FREE #<CONS 0 13573>
 "00000000000000000011010100000110", -- 13573 FREE #<CONS 0 13574>
 "00000000000000000011010100000111", -- 13574 FREE #<CONS 0 13575>
 "00000000000000000011010100001000", -- 13575 FREE #<CONS 0 13576>
 "00000000000000000011010100001001", -- 13576 FREE #<CONS 0 13577>
 "00000000000000000011010100001010", -- 13577 FREE #<CONS 0 13578>
 "00000000000000000011010100001011", -- 13578 FREE #<CONS 0 13579>
 "00000000000000000011010100001100", -- 13579 FREE #<CONS 0 13580>
 "00000000000000000011010100001101", -- 13580 FREE #<CONS 0 13581>
 "00000000000000000011010100001110", -- 13581 FREE #<CONS 0 13582>
 "00000000000000000011010100001111", -- 13582 FREE #<CONS 0 13583>
 "00000000000000000011010100010000", -- 13583 FREE #<CONS 0 13584>
 "00000000000000000011010100010001", -- 13584 FREE #<CONS 0 13585>
 "00000000000000000011010100010010", -- 13585 FREE #<CONS 0 13586>
 "00000000000000000011010100010011", -- 13586 FREE #<CONS 0 13587>
 "00000000000000000011010100010100", -- 13587 FREE #<CONS 0 13588>
 "00000000000000000011010100010101", -- 13588 FREE #<CONS 0 13589>
 "00000000000000000011010100010110", -- 13589 FREE #<CONS 0 13590>
 "00000000000000000011010100010111", -- 13590 FREE #<CONS 0 13591>
 "00000000000000000011010100011000", -- 13591 FREE #<CONS 0 13592>
 "00000000000000000011010100011001", -- 13592 FREE #<CONS 0 13593>
 "00000000000000000011010100011010", -- 13593 FREE #<CONS 0 13594>
 "00000000000000000011010100011011", -- 13594 FREE #<CONS 0 13595>
 "00000000000000000011010100011100", -- 13595 FREE #<CONS 0 13596>
 "00000000000000000011010100011101", -- 13596 FREE #<CONS 0 13597>
 "00000000000000000011010100011110", -- 13597 FREE #<CONS 0 13598>
 "00000000000000000011010100011111", -- 13598 FREE #<CONS 0 13599>
 "00000000000000000011010100100000", -- 13599 FREE #<CONS 0 13600>
 "00000000000000000011010100100001", -- 13600 FREE #<CONS 0 13601>
 "00000000000000000011010100100010", -- 13601 FREE #<CONS 0 13602>
 "00000000000000000011010100100011", -- 13602 FREE #<CONS 0 13603>
 "00000000000000000011010100100100", -- 13603 FREE #<CONS 0 13604>
 "00000000000000000011010100100101", -- 13604 FREE #<CONS 0 13605>
 "00000000000000000011010100100110", -- 13605 FREE #<CONS 0 13606>
 "00000000000000000011010100100111", -- 13606 FREE #<CONS 0 13607>
 "00000000000000000011010100101000", -- 13607 FREE #<CONS 0 13608>
 "00000000000000000011010100101001", -- 13608 FREE #<CONS 0 13609>
 "00000000000000000011010100101010", -- 13609 FREE #<CONS 0 13610>
 "00000000000000000011010100101011", -- 13610 FREE #<CONS 0 13611>
 "00000000000000000011010100101100", -- 13611 FREE #<CONS 0 13612>
 "00000000000000000011010100101101", -- 13612 FREE #<CONS 0 13613>
 "00000000000000000011010100101110", -- 13613 FREE #<CONS 0 13614>
 "00000000000000000011010100101111", -- 13614 FREE #<CONS 0 13615>
 "00000000000000000011010100110000", -- 13615 FREE #<CONS 0 13616>
 "00000000000000000011010100110001", -- 13616 FREE #<CONS 0 13617>
 "00000000000000000011010100110010", -- 13617 FREE #<CONS 0 13618>
 "00000000000000000011010100110011", -- 13618 FREE #<CONS 0 13619>
 "00000000000000000011010100110100", -- 13619 FREE #<CONS 0 13620>
 "00000000000000000011010100110101", -- 13620 FREE #<CONS 0 13621>
 "00000000000000000011010100110110", -- 13621 FREE #<CONS 0 13622>
 "00000000000000000011010100110111", -- 13622 FREE #<CONS 0 13623>
 "00000000000000000011010100111000", -- 13623 FREE #<CONS 0 13624>
 "00000000000000000011010100111001", -- 13624 FREE #<CONS 0 13625>
 "00000000000000000011010100111010", -- 13625 FREE #<CONS 0 13626>
 "00000000000000000011010100111011", -- 13626 FREE #<CONS 0 13627>
 "00000000000000000011010100111100", -- 13627 FREE #<CONS 0 13628>
 "00000000000000000011010100111101", -- 13628 FREE #<CONS 0 13629>
 "00000000000000000011010100111110", -- 13629 FREE #<CONS 0 13630>
 "00000000000000000011010100111111", -- 13630 FREE #<CONS 0 13631>
 "00000000000000000011010101000000", -- 13631 FREE #<CONS 0 13632>
 "00000000000000000011010101000001", -- 13632 FREE #<CONS 0 13633>
 "00000000000000000011010101000010", -- 13633 FREE #<CONS 0 13634>
 "00000000000000000011010101000011", -- 13634 FREE #<CONS 0 13635>
 "00000000000000000011010101000100", -- 13635 FREE #<CONS 0 13636>
 "00000000000000000011010101000101", -- 13636 FREE #<CONS 0 13637>
 "00000000000000000011010101000110", -- 13637 FREE #<CONS 0 13638>
 "00000000000000000011010101000111", -- 13638 FREE #<CONS 0 13639>
 "00000000000000000011010101001000", -- 13639 FREE #<CONS 0 13640>
 "00000000000000000011010101001001", -- 13640 FREE #<CONS 0 13641>
 "00000000000000000011010101001010", -- 13641 FREE #<CONS 0 13642>
 "00000000000000000011010101001011", -- 13642 FREE #<CONS 0 13643>
 "00000000000000000011010101001100", -- 13643 FREE #<CONS 0 13644>
 "00000000000000000011010101001101", -- 13644 FREE #<CONS 0 13645>
 "00000000000000000011010101001110", -- 13645 FREE #<CONS 0 13646>
 "00000000000000000011010101001111", -- 13646 FREE #<CONS 0 13647>
 "00000000000000000011010101010000", -- 13647 FREE #<CONS 0 13648>
 "00000000000000000011010101010001", -- 13648 FREE #<CONS 0 13649>
 "00000000000000000011010101010010", -- 13649 FREE #<CONS 0 13650>
 "00000000000000000011010101010011", -- 13650 FREE #<CONS 0 13651>
 "00000000000000000011010101010100", -- 13651 FREE #<CONS 0 13652>
 "00000000000000000011010101010101", -- 13652 FREE #<CONS 0 13653>
 "00000000000000000011010101010110", -- 13653 FREE #<CONS 0 13654>
 "00000000000000000011010101010111", -- 13654 FREE #<CONS 0 13655>
 "00000000000000000011010101011000", -- 13655 FREE #<CONS 0 13656>
 "00000000000000000011010101011001", -- 13656 FREE #<CONS 0 13657>
 "00000000000000000011010101011010", -- 13657 FREE #<CONS 0 13658>
 "00000000000000000011010101011011", -- 13658 FREE #<CONS 0 13659>
 "00000000000000000011010101011100", -- 13659 FREE #<CONS 0 13660>
 "00000000000000000011010101011101", -- 13660 FREE #<CONS 0 13661>
 "00000000000000000011010101011110", -- 13661 FREE #<CONS 0 13662>
 "00000000000000000011010101011111", -- 13662 FREE #<CONS 0 13663>
 "00000000000000000011010101100000", -- 13663 FREE #<CONS 0 13664>
 "00000000000000000011010101100001", -- 13664 FREE #<CONS 0 13665>
 "00000000000000000011010101100010", -- 13665 FREE #<CONS 0 13666>
 "00000000000000000011010101100011", -- 13666 FREE #<CONS 0 13667>
 "00000000000000000011010101100100", -- 13667 FREE #<CONS 0 13668>
 "00000000000000000011010101100101", -- 13668 FREE #<CONS 0 13669>
 "00000000000000000011010101100110", -- 13669 FREE #<CONS 0 13670>
 "00000000000000000011010101100111", -- 13670 FREE #<CONS 0 13671>
 "00000000000000000011010101101000", -- 13671 FREE #<CONS 0 13672>
 "00000000000000000011010101101001", -- 13672 FREE #<CONS 0 13673>
 "00000000000000000011010101101010", -- 13673 FREE #<CONS 0 13674>
 "00000000000000000011010101101011", -- 13674 FREE #<CONS 0 13675>
 "00000000000000000011010101101100", -- 13675 FREE #<CONS 0 13676>
 "00000000000000000011010101101101", -- 13676 FREE #<CONS 0 13677>
 "00000000000000000011010101101110", -- 13677 FREE #<CONS 0 13678>
 "00000000000000000011010101101111", -- 13678 FREE #<CONS 0 13679>
 "00000000000000000011010101110000", -- 13679 FREE #<CONS 0 13680>
 "00000000000000000011010101110001", -- 13680 FREE #<CONS 0 13681>
 "00000000000000000011010101110010", -- 13681 FREE #<CONS 0 13682>
 "00000000000000000011010101110011", -- 13682 FREE #<CONS 0 13683>
 "00000000000000000011010101110100", -- 13683 FREE #<CONS 0 13684>
 "00000000000000000011010101110101", -- 13684 FREE #<CONS 0 13685>
 "00000000000000000011010101110110", -- 13685 FREE #<CONS 0 13686>
 "00000000000000000011010101110111", -- 13686 FREE #<CONS 0 13687>
 "00000000000000000011010101111000", -- 13687 FREE #<CONS 0 13688>
 "00000000000000000011010101111001", -- 13688 FREE #<CONS 0 13689>
 "00000000000000000011010101111010", -- 13689 FREE #<CONS 0 13690>
 "00000000000000000011010101111011", -- 13690 FREE #<CONS 0 13691>
 "00000000000000000011010101111100", -- 13691 FREE #<CONS 0 13692>
 "00000000000000000011010101111101", -- 13692 FREE #<CONS 0 13693>
 "00000000000000000011010101111110", -- 13693 FREE #<CONS 0 13694>
 "00000000000000000011010101111111", -- 13694 FREE #<CONS 0 13695>
 "00000000000000000011010110000000", -- 13695 FREE #<CONS 0 13696>
 "00000000000000000011010110000001", -- 13696 FREE #<CONS 0 13697>
 "00000000000000000011010110000010", -- 13697 FREE #<CONS 0 13698>
 "00000000000000000011010110000011", -- 13698 FREE #<CONS 0 13699>
 "00000000000000000011010110000100", -- 13699 FREE #<CONS 0 13700>
 "00000000000000000011010110000101", -- 13700 FREE #<CONS 0 13701>
 "00000000000000000011010110000110", -- 13701 FREE #<CONS 0 13702>
 "00000000000000000011010110000111", -- 13702 FREE #<CONS 0 13703>
 "00000000000000000011010110001000", -- 13703 FREE #<CONS 0 13704>
 "00000000000000000011010110001001", -- 13704 FREE #<CONS 0 13705>
 "00000000000000000011010110001010", -- 13705 FREE #<CONS 0 13706>
 "00000000000000000011010110001011", -- 13706 FREE #<CONS 0 13707>
 "00000000000000000011010110001100", -- 13707 FREE #<CONS 0 13708>
 "00000000000000000011010110001101", -- 13708 FREE #<CONS 0 13709>
 "00000000000000000011010110001110", -- 13709 FREE #<CONS 0 13710>
 "00000000000000000011010110001111", -- 13710 FREE #<CONS 0 13711>
 "00000000000000000011010110010000", -- 13711 FREE #<CONS 0 13712>
 "00000000000000000011010110010001", -- 13712 FREE #<CONS 0 13713>
 "00000000000000000011010110010010", -- 13713 FREE #<CONS 0 13714>
 "00000000000000000011010110010011", -- 13714 FREE #<CONS 0 13715>
 "00000000000000000011010110010100", -- 13715 FREE #<CONS 0 13716>
 "00000000000000000011010110010101", -- 13716 FREE #<CONS 0 13717>
 "00000000000000000011010110010110", -- 13717 FREE #<CONS 0 13718>
 "00000000000000000011010110010111", -- 13718 FREE #<CONS 0 13719>
 "00000000000000000011010110011000", -- 13719 FREE #<CONS 0 13720>
 "00000000000000000011010110011001", -- 13720 FREE #<CONS 0 13721>
 "00000000000000000011010110011010", -- 13721 FREE #<CONS 0 13722>
 "00000000000000000011010110011011", -- 13722 FREE #<CONS 0 13723>
 "00000000000000000011010110011100", -- 13723 FREE #<CONS 0 13724>
 "00000000000000000011010110011101", -- 13724 FREE #<CONS 0 13725>
 "00000000000000000011010110011110", -- 13725 FREE #<CONS 0 13726>
 "00000000000000000011010110011111", -- 13726 FREE #<CONS 0 13727>
 "00000000000000000011010110100000", -- 13727 FREE #<CONS 0 13728>
 "00000000000000000011010110100001", -- 13728 FREE #<CONS 0 13729>
 "00000000000000000011010110100010", -- 13729 FREE #<CONS 0 13730>
 "00000000000000000011010110100011", -- 13730 FREE #<CONS 0 13731>
 "00000000000000000011010110100100", -- 13731 FREE #<CONS 0 13732>
 "00000000000000000011010110100101", -- 13732 FREE #<CONS 0 13733>
 "00000000000000000011010110100110", -- 13733 FREE #<CONS 0 13734>
 "00000000000000000011010110100111", -- 13734 FREE #<CONS 0 13735>
 "00000000000000000011010110101000", -- 13735 FREE #<CONS 0 13736>
 "00000000000000000011010110101001", -- 13736 FREE #<CONS 0 13737>
 "00000000000000000011010110101010", -- 13737 FREE #<CONS 0 13738>
 "00000000000000000011010110101011", -- 13738 FREE #<CONS 0 13739>
 "00000000000000000011010110101100", -- 13739 FREE #<CONS 0 13740>
 "00000000000000000011010110101101", -- 13740 FREE #<CONS 0 13741>
 "00000000000000000011010110101110", -- 13741 FREE #<CONS 0 13742>
 "00000000000000000011010110101111", -- 13742 FREE #<CONS 0 13743>
 "00000000000000000011010110110000", -- 13743 FREE #<CONS 0 13744>
 "00000000000000000011010110110001", -- 13744 FREE #<CONS 0 13745>
 "00000000000000000011010110110010", -- 13745 FREE #<CONS 0 13746>
 "00000000000000000011010110110011", -- 13746 FREE #<CONS 0 13747>
 "00000000000000000011010110110100", -- 13747 FREE #<CONS 0 13748>
 "00000000000000000011010110110101", -- 13748 FREE #<CONS 0 13749>
 "00000000000000000011010110110110", -- 13749 FREE #<CONS 0 13750>
 "00000000000000000011010110110111", -- 13750 FREE #<CONS 0 13751>
 "00000000000000000011010110111000", -- 13751 FREE #<CONS 0 13752>
 "00000000000000000011010110111001", -- 13752 FREE #<CONS 0 13753>
 "00000000000000000011010110111010", -- 13753 FREE #<CONS 0 13754>
 "00000000000000000011010110111011", -- 13754 FREE #<CONS 0 13755>
 "00000000000000000011010110111100", -- 13755 FREE #<CONS 0 13756>
 "00000000000000000011010110111101", -- 13756 FREE #<CONS 0 13757>
 "00000000000000000011010110111110", -- 13757 FREE #<CONS 0 13758>
 "00000000000000000011010110111111", -- 13758 FREE #<CONS 0 13759>
 "00000000000000000011010111000000", -- 13759 FREE #<CONS 0 13760>
 "00000000000000000011010111000001", -- 13760 FREE #<CONS 0 13761>
 "00000000000000000011010111000010", -- 13761 FREE #<CONS 0 13762>
 "00000000000000000011010111000011", -- 13762 FREE #<CONS 0 13763>
 "00000000000000000011010111000100", -- 13763 FREE #<CONS 0 13764>
 "00000000000000000011010111000101", -- 13764 FREE #<CONS 0 13765>
 "00000000000000000011010111000110", -- 13765 FREE #<CONS 0 13766>
 "00000000000000000011010111000111", -- 13766 FREE #<CONS 0 13767>
 "00000000000000000011010111001000", -- 13767 FREE #<CONS 0 13768>
 "00000000000000000011010111001001", -- 13768 FREE #<CONS 0 13769>
 "00000000000000000011010111001010", -- 13769 FREE #<CONS 0 13770>
 "00000000000000000011010111001011", -- 13770 FREE #<CONS 0 13771>
 "00000000000000000011010111001100", -- 13771 FREE #<CONS 0 13772>
 "00000000000000000011010111001101", -- 13772 FREE #<CONS 0 13773>
 "00000000000000000011010111001110", -- 13773 FREE #<CONS 0 13774>
 "00000000000000000011010111001111", -- 13774 FREE #<CONS 0 13775>
 "00000000000000000011010111010000", -- 13775 FREE #<CONS 0 13776>
 "00000000000000000011010111010001", -- 13776 FREE #<CONS 0 13777>
 "00000000000000000011010111010010", -- 13777 FREE #<CONS 0 13778>
 "00000000000000000011010111010011", -- 13778 FREE #<CONS 0 13779>
 "00000000000000000011010111010100", -- 13779 FREE #<CONS 0 13780>
 "00000000000000000011010111010101", -- 13780 FREE #<CONS 0 13781>
 "00000000000000000011010111010110", -- 13781 FREE #<CONS 0 13782>
 "00000000000000000011010111010111", -- 13782 FREE #<CONS 0 13783>
 "00000000000000000011010111011000", -- 13783 FREE #<CONS 0 13784>
 "00000000000000000011010111011001", -- 13784 FREE #<CONS 0 13785>
 "00000000000000000011010111011010", -- 13785 FREE #<CONS 0 13786>
 "00000000000000000011010111011011", -- 13786 FREE #<CONS 0 13787>
 "00000000000000000011010111011100", -- 13787 FREE #<CONS 0 13788>
 "00000000000000000011010111011101", -- 13788 FREE #<CONS 0 13789>
 "00000000000000000011010111011110", -- 13789 FREE #<CONS 0 13790>
 "00000000000000000011010111011111", -- 13790 FREE #<CONS 0 13791>
 "00000000000000000011010111100000", -- 13791 FREE #<CONS 0 13792>
 "00000000000000000011010111100001", -- 13792 FREE #<CONS 0 13793>
 "00000000000000000011010111100010", -- 13793 FREE #<CONS 0 13794>
 "00000000000000000011010111100011", -- 13794 FREE #<CONS 0 13795>
 "00000000000000000011010111100100", -- 13795 FREE #<CONS 0 13796>
 "00000000000000000011010111100101", -- 13796 FREE #<CONS 0 13797>
 "00000000000000000011010111100110", -- 13797 FREE #<CONS 0 13798>
 "00000000000000000011010111100111", -- 13798 FREE #<CONS 0 13799>
 "00000000000000000011010111101000", -- 13799 FREE #<CONS 0 13800>
 "00000000000000000011010111101001", -- 13800 FREE #<CONS 0 13801>
 "00000000000000000011010111101010", -- 13801 FREE #<CONS 0 13802>
 "00000000000000000011010111101011", -- 13802 FREE #<CONS 0 13803>
 "00000000000000000011010111101100", -- 13803 FREE #<CONS 0 13804>
 "00000000000000000011010111101101", -- 13804 FREE #<CONS 0 13805>
 "00000000000000000011010111101110", -- 13805 FREE #<CONS 0 13806>
 "00000000000000000011010111101111", -- 13806 FREE #<CONS 0 13807>
 "00000000000000000011010111110000", -- 13807 FREE #<CONS 0 13808>
 "00000000000000000011010111110001", -- 13808 FREE #<CONS 0 13809>
 "00000000000000000011010111110010", -- 13809 FREE #<CONS 0 13810>
 "00000000000000000011010111110011", -- 13810 FREE #<CONS 0 13811>
 "00000000000000000011010111110100", -- 13811 FREE #<CONS 0 13812>
 "00000000000000000011010111110101", -- 13812 FREE #<CONS 0 13813>
 "00000000000000000011010111110110", -- 13813 FREE #<CONS 0 13814>
 "00000000000000000011010111110111", -- 13814 FREE #<CONS 0 13815>
 "00000000000000000011010111111000", -- 13815 FREE #<CONS 0 13816>
 "00000000000000000011010111111001", -- 13816 FREE #<CONS 0 13817>
 "00000000000000000011010111111010", -- 13817 FREE #<CONS 0 13818>
 "00000000000000000011010111111011", -- 13818 FREE #<CONS 0 13819>
 "00000000000000000011010111111100", -- 13819 FREE #<CONS 0 13820>
 "00000000000000000011010111111101", -- 13820 FREE #<CONS 0 13821>
 "00000000000000000011010111111110", -- 13821 FREE #<CONS 0 13822>
 "00000000000000000011010111111111", -- 13822 FREE #<CONS 0 13823>
 "00000000000000000011011000000000", -- 13823 FREE #<CONS 0 13824>
 "00000000000000000011011000000001", -- 13824 FREE #<CONS 0 13825>
 "00000000000000000011011000000010", -- 13825 FREE #<CONS 0 13826>
 "00000000000000000011011000000011", -- 13826 FREE #<CONS 0 13827>
 "00000000000000000011011000000100", -- 13827 FREE #<CONS 0 13828>
 "00000000000000000011011000000101", -- 13828 FREE #<CONS 0 13829>
 "00000000000000000011011000000110", -- 13829 FREE #<CONS 0 13830>
 "00000000000000000011011000000111", -- 13830 FREE #<CONS 0 13831>
 "00000000000000000011011000001000", -- 13831 FREE #<CONS 0 13832>
 "00000000000000000011011000001001", -- 13832 FREE #<CONS 0 13833>
 "00000000000000000011011000001010", -- 13833 FREE #<CONS 0 13834>
 "00000000000000000011011000001011", -- 13834 FREE #<CONS 0 13835>
 "00000000000000000011011000001100", -- 13835 FREE #<CONS 0 13836>
 "00000000000000000011011000001101", -- 13836 FREE #<CONS 0 13837>
 "00000000000000000011011000001110", -- 13837 FREE #<CONS 0 13838>
 "00000000000000000011011000001111", -- 13838 FREE #<CONS 0 13839>
 "00000000000000000011011000010000", -- 13839 FREE #<CONS 0 13840>
 "00000000000000000011011000010001", -- 13840 FREE #<CONS 0 13841>
 "00000000000000000011011000010010", -- 13841 FREE #<CONS 0 13842>
 "00000000000000000011011000010011", -- 13842 FREE #<CONS 0 13843>
 "00000000000000000011011000010100", -- 13843 FREE #<CONS 0 13844>
 "00000000000000000011011000010101", -- 13844 FREE #<CONS 0 13845>
 "00000000000000000011011000010110", -- 13845 FREE #<CONS 0 13846>
 "00000000000000000011011000010111", -- 13846 FREE #<CONS 0 13847>
 "00000000000000000011011000011000", -- 13847 FREE #<CONS 0 13848>
 "00000000000000000011011000011001", -- 13848 FREE #<CONS 0 13849>
 "00000000000000000011011000011010", -- 13849 FREE #<CONS 0 13850>
 "00000000000000000011011000011011", -- 13850 FREE #<CONS 0 13851>
 "00000000000000000011011000011100", -- 13851 FREE #<CONS 0 13852>
 "00000000000000000011011000011101", -- 13852 FREE #<CONS 0 13853>
 "00000000000000000011011000011110", -- 13853 FREE #<CONS 0 13854>
 "00000000000000000011011000011111", -- 13854 FREE #<CONS 0 13855>
 "00000000000000000011011000100000", -- 13855 FREE #<CONS 0 13856>
 "00000000000000000011011000100001", -- 13856 FREE #<CONS 0 13857>
 "00000000000000000011011000100010", -- 13857 FREE #<CONS 0 13858>
 "00000000000000000011011000100011", -- 13858 FREE #<CONS 0 13859>
 "00000000000000000011011000100100", -- 13859 FREE #<CONS 0 13860>
 "00000000000000000011011000100101", -- 13860 FREE #<CONS 0 13861>
 "00000000000000000011011000100110", -- 13861 FREE #<CONS 0 13862>
 "00000000000000000011011000100111", -- 13862 FREE #<CONS 0 13863>
 "00000000000000000011011000101000", -- 13863 FREE #<CONS 0 13864>
 "00000000000000000011011000101001", -- 13864 FREE #<CONS 0 13865>
 "00000000000000000011011000101010", -- 13865 FREE #<CONS 0 13866>
 "00000000000000000011011000101011", -- 13866 FREE #<CONS 0 13867>
 "00000000000000000011011000101100", -- 13867 FREE #<CONS 0 13868>
 "00000000000000000011011000101101", -- 13868 FREE #<CONS 0 13869>
 "00000000000000000011011000101110", -- 13869 FREE #<CONS 0 13870>
 "00000000000000000011011000101111", -- 13870 FREE #<CONS 0 13871>
 "00000000000000000011011000110000", -- 13871 FREE #<CONS 0 13872>
 "00000000000000000011011000110001", -- 13872 FREE #<CONS 0 13873>
 "00000000000000000011011000110010", -- 13873 FREE #<CONS 0 13874>
 "00000000000000000011011000110011", -- 13874 FREE #<CONS 0 13875>
 "00000000000000000011011000110100", -- 13875 FREE #<CONS 0 13876>
 "00000000000000000011011000110101", -- 13876 FREE #<CONS 0 13877>
 "00000000000000000011011000110110", -- 13877 FREE #<CONS 0 13878>
 "00000000000000000011011000110111", -- 13878 FREE #<CONS 0 13879>
 "00000000000000000011011000111000", -- 13879 FREE #<CONS 0 13880>
 "00000000000000000011011000111001", -- 13880 FREE #<CONS 0 13881>
 "00000000000000000011011000111010", -- 13881 FREE #<CONS 0 13882>
 "00000000000000000011011000111011", -- 13882 FREE #<CONS 0 13883>
 "00000000000000000011011000111100", -- 13883 FREE #<CONS 0 13884>
 "00000000000000000011011000111101", -- 13884 FREE #<CONS 0 13885>
 "00000000000000000011011000111110", -- 13885 FREE #<CONS 0 13886>
 "00000000000000000011011000111111", -- 13886 FREE #<CONS 0 13887>
 "00000000000000000011011001000000", -- 13887 FREE #<CONS 0 13888>
 "00000000000000000011011001000001", -- 13888 FREE #<CONS 0 13889>
 "00000000000000000011011001000010", -- 13889 FREE #<CONS 0 13890>
 "00000000000000000011011001000011", -- 13890 FREE #<CONS 0 13891>
 "00000000000000000011011001000100", -- 13891 FREE #<CONS 0 13892>
 "00000000000000000011011001000101", -- 13892 FREE #<CONS 0 13893>
 "00000000000000000011011001000110", -- 13893 FREE #<CONS 0 13894>
 "00000000000000000011011001000111", -- 13894 FREE #<CONS 0 13895>
 "00000000000000000011011001001000", -- 13895 FREE #<CONS 0 13896>
 "00000000000000000011011001001001", -- 13896 FREE #<CONS 0 13897>
 "00000000000000000011011001001010", -- 13897 FREE #<CONS 0 13898>
 "00000000000000000011011001001011", -- 13898 FREE #<CONS 0 13899>
 "00000000000000000011011001001100", -- 13899 FREE #<CONS 0 13900>
 "00000000000000000011011001001101", -- 13900 FREE #<CONS 0 13901>
 "00000000000000000011011001001110", -- 13901 FREE #<CONS 0 13902>
 "00000000000000000011011001001111", -- 13902 FREE #<CONS 0 13903>
 "00000000000000000011011001010000", -- 13903 FREE #<CONS 0 13904>
 "00000000000000000011011001010001", -- 13904 FREE #<CONS 0 13905>
 "00000000000000000011011001010010", -- 13905 FREE #<CONS 0 13906>
 "00000000000000000011011001010011", -- 13906 FREE #<CONS 0 13907>
 "00000000000000000011011001010100", -- 13907 FREE #<CONS 0 13908>
 "00000000000000000011011001010101", -- 13908 FREE #<CONS 0 13909>
 "00000000000000000011011001010110", -- 13909 FREE #<CONS 0 13910>
 "00000000000000000011011001010111", -- 13910 FREE #<CONS 0 13911>
 "00000000000000000011011001011000", -- 13911 FREE #<CONS 0 13912>
 "00000000000000000011011001011001", -- 13912 FREE #<CONS 0 13913>
 "00000000000000000011011001011010", -- 13913 FREE #<CONS 0 13914>
 "00000000000000000011011001011011", -- 13914 FREE #<CONS 0 13915>
 "00000000000000000011011001011100", -- 13915 FREE #<CONS 0 13916>
 "00000000000000000011011001011101", -- 13916 FREE #<CONS 0 13917>
 "00000000000000000011011001011110", -- 13917 FREE #<CONS 0 13918>
 "00000000000000000011011001011111", -- 13918 FREE #<CONS 0 13919>
 "00000000000000000011011001100000", -- 13919 FREE #<CONS 0 13920>
 "00000000000000000011011001100001", -- 13920 FREE #<CONS 0 13921>
 "00000000000000000011011001100010", -- 13921 FREE #<CONS 0 13922>
 "00000000000000000011011001100011", -- 13922 FREE #<CONS 0 13923>
 "00000000000000000011011001100100", -- 13923 FREE #<CONS 0 13924>
 "00000000000000000011011001100101", -- 13924 FREE #<CONS 0 13925>
 "00000000000000000011011001100110", -- 13925 FREE #<CONS 0 13926>
 "00000000000000000011011001100111", -- 13926 FREE #<CONS 0 13927>
 "00000000000000000011011001101000", -- 13927 FREE #<CONS 0 13928>
 "00000000000000000011011001101001", -- 13928 FREE #<CONS 0 13929>
 "00000000000000000011011001101010", -- 13929 FREE #<CONS 0 13930>
 "00000000000000000011011001101011", -- 13930 FREE #<CONS 0 13931>
 "00000000000000000011011001101100", -- 13931 FREE #<CONS 0 13932>
 "00000000000000000011011001101101", -- 13932 FREE #<CONS 0 13933>
 "00000000000000000011011001101110", -- 13933 FREE #<CONS 0 13934>
 "00000000000000000011011001101111", -- 13934 FREE #<CONS 0 13935>
 "00000000000000000011011001110000", -- 13935 FREE #<CONS 0 13936>
 "00000000000000000011011001110001", -- 13936 FREE #<CONS 0 13937>
 "00000000000000000011011001110010", -- 13937 FREE #<CONS 0 13938>
 "00000000000000000011011001110011", -- 13938 FREE #<CONS 0 13939>
 "00000000000000000011011001110100", -- 13939 FREE #<CONS 0 13940>
 "00000000000000000011011001110101", -- 13940 FREE #<CONS 0 13941>
 "00000000000000000011011001110110", -- 13941 FREE #<CONS 0 13942>
 "00000000000000000011011001110111", -- 13942 FREE #<CONS 0 13943>
 "00000000000000000011011001111000", -- 13943 FREE #<CONS 0 13944>
 "00000000000000000011011001111001", -- 13944 FREE #<CONS 0 13945>
 "00000000000000000011011001111010", -- 13945 FREE #<CONS 0 13946>
 "00000000000000000011011001111011", -- 13946 FREE #<CONS 0 13947>
 "00000000000000000011011001111100", -- 13947 FREE #<CONS 0 13948>
 "00000000000000000011011001111101", -- 13948 FREE #<CONS 0 13949>
 "00000000000000000011011001111110", -- 13949 FREE #<CONS 0 13950>
 "00000000000000000011011001111111", -- 13950 FREE #<CONS 0 13951>
 "00000000000000000011011010000000", -- 13951 FREE #<CONS 0 13952>
 "00000000000000000011011010000001", -- 13952 FREE #<CONS 0 13953>
 "00000000000000000011011010000010", -- 13953 FREE #<CONS 0 13954>
 "00000000000000000011011010000011", -- 13954 FREE #<CONS 0 13955>
 "00000000000000000011011010000100", -- 13955 FREE #<CONS 0 13956>
 "00000000000000000011011010000101", -- 13956 FREE #<CONS 0 13957>
 "00000000000000000011011010000110", -- 13957 FREE #<CONS 0 13958>
 "00000000000000000011011010000111", -- 13958 FREE #<CONS 0 13959>
 "00000000000000000011011010001000", -- 13959 FREE #<CONS 0 13960>
 "00000000000000000011011010001001", -- 13960 FREE #<CONS 0 13961>
 "00000000000000000011011010001010", -- 13961 FREE #<CONS 0 13962>
 "00000000000000000011011010001011", -- 13962 FREE #<CONS 0 13963>
 "00000000000000000011011010001100", -- 13963 FREE #<CONS 0 13964>
 "00000000000000000011011010001101", -- 13964 FREE #<CONS 0 13965>
 "00000000000000000011011010001110", -- 13965 FREE #<CONS 0 13966>
 "00000000000000000011011010001111", -- 13966 FREE #<CONS 0 13967>
 "00000000000000000011011010010000", -- 13967 FREE #<CONS 0 13968>
 "00000000000000000011011010010001", -- 13968 FREE #<CONS 0 13969>
 "00000000000000000011011010010010", -- 13969 FREE #<CONS 0 13970>
 "00000000000000000011011010010011", -- 13970 FREE #<CONS 0 13971>
 "00000000000000000011011010010100", -- 13971 FREE #<CONS 0 13972>
 "00000000000000000011011010010101", -- 13972 FREE #<CONS 0 13973>
 "00000000000000000011011010010110", -- 13973 FREE #<CONS 0 13974>
 "00000000000000000011011010010111", -- 13974 FREE #<CONS 0 13975>
 "00000000000000000011011010011000", -- 13975 FREE #<CONS 0 13976>
 "00000000000000000011011010011001", -- 13976 FREE #<CONS 0 13977>
 "00000000000000000011011010011010", -- 13977 FREE #<CONS 0 13978>
 "00000000000000000011011010011011", -- 13978 FREE #<CONS 0 13979>
 "00000000000000000011011010011100", -- 13979 FREE #<CONS 0 13980>
 "00000000000000000011011010011101", -- 13980 FREE #<CONS 0 13981>
 "00000000000000000011011010011110", -- 13981 FREE #<CONS 0 13982>
 "00000000000000000011011010011111", -- 13982 FREE #<CONS 0 13983>
 "00000000000000000011011010100000", -- 13983 FREE #<CONS 0 13984>
 "00000000000000000011011010100001", -- 13984 FREE #<CONS 0 13985>
 "00000000000000000011011010100010", -- 13985 FREE #<CONS 0 13986>
 "00000000000000000011011010100011", -- 13986 FREE #<CONS 0 13987>
 "00000000000000000011011010100100", -- 13987 FREE #<CONS 0 13988>
 "00000000000000000011011010100101", -- 13988 FREE #<CONS 0 13989>
 "00000000000000000011011010100110", -- 13989 FREE #<CONS 0 13990>
 "00000000000000000011011010100111", -- 13990 FREE #<CONS 0 13991>
 "00000000000000000011011010101000", -- 13991 FREE #<CONS 0 13992>
 "00000000000000000011011010101001", -- 13992 FREE #<CONS 0 13993>
 "00000000000000000011011010101010", -- 13993 FREE #<CONS 0 13994>
 "00000000000000000011011010101011", -- 13994 FREE #<CONS 0 13995>
 "00000000000000000011011010101100", -- 13995 FREE #<CONS 0 13996>
 "00000000000000000011011010101101", -- 13996 FREE #<CONS 0 13997>
 "00000000000000000011011010101110", -- 13997 FREE #<CONS 0 13998>
 "00000000000000000011011010101111", -- 13998 FREE #<CONS 0 13999>
 "00000000000000000011011010110000", -- 13999 FREE #<CONS 0 14000>
 "00000000000000000011011010110001", -- 14000 FREE #<CONS 0 14001>
 "00000000000000000011011010110010", -- 14001 FREE #<CONS 0 14002>
 "00000000000000000011011010110011", -- 14002 FREE #<CONS 0 14003>
 "00000000000000000011011010110100", -- 14003 FREE #<CONS 0 14004>
 "00000000000000000011011010110101", -- 14004 FREE #<CONS 0 14005>
 "00000000000000000011011010110110", -- 14005 FREE #<CONS 0 14006>
 "00000000000000000011011010110111", -- 14006 FREE #<CONS 0 14007>
 "00000000000000000011011010111000", -- 14007 FREE #<CONS 0 14008>
 "00000000000000000011011010111001", -- 14008 FREE #<CONS 0 14009>
 "00000000000000000011011010111010", -- 14009 FREE #<CONS 0 14010>
 "00000000000000000011011010111011", -- 14010 FREE #<CONS 0 14011>
 "00000000000000000011011010111100", -- 14011 FREE #<CONS 0 14012>
 "00000000000000000011011010111101", -- 14012 FREE #<CONS 0 14013>
 "00000000000000000011011010111110", -- 14013 FREE #<CONS 0 14014>
 "00000000000000000011011010111111", -- 14014 FREE #<CONS 0 14015>
 "00000000000000000011011011000000", -- 14015 FREE #<CONS 0 14016>
 "00000000000000000011011011000001", -- 14016 FREE #<CONS 0 14017>
 "00000000000000000011011011000010", -- 14017 FREE #<CONS 0 14018>
 "00000000000000000011011011000011", -- 14018 FREE #<CONS 0 14019>
 "00000000000000000011011011000100", -- 14019 FREE #<CONS 0 14020>
 "00000000000000000011011011000101", -- 14020 FREE #<CONS 0 14021>
 "00000000000000000011011011000110", -- 14021 FREE #<CONS 0 14022>
 "00000000000000000011011011000111", -- 14022 FREE #<CONS 0 14023>
 "00000000000000000011011011001000", -- 14023 FREE #<CONS 0 14024>
 "00000000000000000011011011001001", -- 14024 FREE #<CONS 0 14025>
 "00000000000000000011011011001010", -- 14025 FREE #<CONS 0 14026>
 "00000000000000000011011011001011", -- 14026 FREE #<CONS 0 14027>
 "00000000000000000011011011001100", -- 14027 FREE #<CONS 0 14028>
 "00000000000000000011011011001101", -- 14028 FREE #<CONS 0 14029>
 "00000000000000000011011011001110", -- 14029 FREE #<CONS 0 14030>
 "00000000000000000011011011001111", -- 14030 FREE #<CONS 0 14031>
 "00000000000000000011011011010000", -- 14031 FREE #<CONS 0 14032>
 "00000000000000000011011011010001", -- 14032 FREE #<CONS 0 14033>
 "00000000000000000011011011010010", -- 14033 FREE #<CONS 0 14034>
 "00000000000000000011011011010011", -- 14034 FREE #<CONS 0 14035>
 "00000000000000000011011011010100", -- 14035 FREE #<CONS 0 14036>
 "00000000000000000011011011010101", -- 14036 FREE #<CONS 0 14037>
 "00000000000000000011011011010110", -- 14037 FREE #<CONS 0 14038>
 "00000000000000000011011011010111", -- 14038 FREE #<CONS 0 14039>
 "00000000000000000011011011011000", -- 14039 FREE #<CONS 0 14040>
 "00000000000000000011011011011001", -- 14040 FREE #<CONS 0 14041>
 "00000000000000000011011011011010", -- 14041 FREE #<CONS 0 14042>
 "00000000000000000011011011011011", -- 14042 FREE #<CONS 0 14043>
 "00000000000000000011011011011100", -- 14043 FREE #<CONS 0 14044>
 "00000000000000000011011011011101", -- 14044 FREE #<CONS 0 14045>
 "00000000000000000011011011011110", -- 14045 FREE #<CONS 0 14046>
 "00000000000000000011011011011111", -- 14046 FREE #<CONS 0 14047>
 "00000000000000000011011011100000", -- 14047 FREE #<CONS 0 14048>
 "00000000000000000011011011100001", -- 14048 FREE #<CONS 0 14049>
 "00000000000000000011011011100010", -- 14049 FREE #<CONS 0 14050>
 "00000000000000000011011011100011", -- 14050 FREE #<CONS 0 14051>
 "00000000000000000011011011100100", -- 14051 FREE #<CONS 0 14052>
 "00000000000000000011011011100101", -- 14052 FREE #<CONS 0 14053>
 "00000000000000000011011011100110", -- 14053 FREE #<CONS 0 14054>
 "00000000000000000011011011100111", -- 14054 FREE #<CONS 0 14055>
 "00000000000000000011011011101000", -- 14055 FREE #<CONS 0 14056>
 "00000000000000000011011011101001", -- 14056 FREE #<CONS 0 14057>
 "00000000000000000011011011101010", -- 14057 FREE #<CONS 0 14058>
 "00000000000000000011011011101011", -- 14058 FREE #<CONS 0 14059>
 "00000000000000000011011011101100", -- 14059 FREE #<CONS 0 14060>
 "00000000000000000011011011101101", -- 14060 FREE #<CONS 0 14061>
 "00000000000000000011011011101110", -- 14061 FREE #<CONS 0 14062>
 "00000000000000000011011011101111", -- 14062 FREE #<CONS 0 14063>
 "00000000000000000011011011110000", -- 14063 FREE #<CONS 0 14064>
 "00000000000000000011011011110001", -- 14064 FREE #<CONS 0 14065>
 "00000000000000000011011011110010", -- 14065 FREE #<CONS 0 14066>
 "00000000000000000011011011110011", -- 14066 FREE #<CONS 0 14067>
 "00000000000000000011011011110100", -- 14067 FREE #<CONS 0 14068>
 "00000000000000000011011011110101", -- 14068 FREE #<CONS 0 14069>
 "00000000000000000011011011110110", -- 14069 FREE #<CONS 0 14070>
 "00000000000000000011011011110111", -- 14070 FREE #<CONS 0 14071>
 "00000000000000000011011011111000", -- 14071 FREE #<CONS 0 14072>
 "00000000000000000011011011111001", -- 14072 FREE #<CONS 0 14073>
 "00000000000000000011011011111010", -- 14073 FREE #<CONS 0 14074>
 "00000000000000000011011011111011", -- 14074 FREE #<CONS 0 14075>
 "00000000000000000011011011111100", -- 14075 FREE #<CONS 0 14076>
 "00000000000000000011011011111101", -- 14076 FREE #<CONS 0 14077>
 "00000000000000000011011011111110", -- 14077 FREE #<CONS 0 14078>
 "00000000000000000011011011111111", -- 14078 FREE #<CONS 0 14079>
 "00000000000000000011011100000000", -- 14079 FREE #<CONS 0 14080>
 "00000000000000000011011100000001", -- 14080 FREE #<CONS 0 14081>
 "00000000000000000011011100000010", -- 14081 FREE #<CONS 0 14082>
 "00000000000000000011011100000011", -- 14082 FREE #<CONS 0 14083>
 "00000000000000000011011100000100", -- 14083 FREE #<CONS 0 14084>
 "00000000000000000011011100000101", -- 14084 FREE #<CONS 0 14085>
 "00000000000000000011011100000110", -- 14085 FREE #<CONS 0 14086>
 "00000000000000000011011100000111", -- 14086 FREE #<CONS 0 14087>
 "00000000000000000011011100001000", -- 14087 FREE #<CONS 0 14088>
 "00000000000000000011011100001001", -- 14088 FREE #<CONS 0 14089>
 "00000000000000000011011100001010", -- 14089 FREE #<CONS 0 14090>
 "00000000000000000011011100001011", -- 14090 FREE #<CONS 0 14091>
 "00000000000000000011011100001100", -- 14091 FREE #<CONS 0 14092>
 "00000000000000000011011100001101", -- 14092 FREE #<CONS 0 14093>
 "00000000000000000011011100001110", -- 14093 FREE #<CONS 0 14094>
 "00000000000000000011011100001111", -- 14094 FREE #<CONS 0 14095>
 "00000000000000000011011100010000", -- 14095 FREE #<CONS 0 14096>
 "00000000000000000011011100010001", -- 14096 FREE #<CONS 0 14097>
 "00000000000000000011011100010010", -- 14097 FREE #<CONS 0 14098>
 "00000000000000000011011100010011", -- 14098 FREE #<CONS 0 14099>
 "00000000000000000011011100010100", -- 14099 FREE #<CONS 0 14100>
 "00000000000000000011011100010101", -- 14100 FREE #<CONS 0 14101>
 "00000000000000000011011100010110", -- 14101 FREE #<CONS 0 14102>
 "00000000000000000011011100010111", -- 14102 FREE #<CONS 0 14103>
 "00000000000000000011011100011000", -- 14103 FREE #<CONS 0 14104>
 "00000000000000000011011100011001", -- 14104 FREE #<CONS 0 14105>
 "00000000000000000011011100011010", -- 14105 FREE #<CONS 0 14106>
 "00000000000000000011011100011011", -- 14106 FREE #<CONS 0 14107>
 "00000000000000000011011100011100", -- 14107 FREE #<CONS 0 14108>
 "00000000000000000011011100011101", -- 14108 FREE #<CONS 0 14109>
 "00000000000000000011011100011110", -- 14109 FREE #<CONS 0 14110>
 "00000000000000000011011100011111", -- 14110 FREE #<CONS 0 14111>
 "00000000000000000011011100100000", -- 14111 FREE #<CONS 0 14112>
 "00000000000000000011011100100001", -- 14112 FREE #<CONS 0 14113>
 "00000000000000000011011100100010", -- 14113 FREE #<CONS 0 14114>
 "00000000000000000011011100100011", -- 14114 FREE #<CONS 0 14115>
 "00000000000000000011011100100100", -- 14115 FREE #<CONS 0 14116>
 "00000000000000000011011100100101", -- 14116 FREE #<CONS 0 14117>
 "00000000000000000011011100100110", -- 14117 FREE #<CONS 0 14118>
 "00000000000000000011011100100111", -- 14118 FREE #<CONS 0 14119>
 "00000000000000000011011100101000", -- 14119 FREE #<CONS 0 14120>
 "00000000000000000011011100101001", -- 14120 FREE #<CONS 0 14121>
 "00000000000000000011011100101010", -- 14121 FREE #<CONS 0 14122>
 "00000000000000000011011100101011", -- 14122 FREE #<CONS 0 14123>
 "00000000000000000011011100101100", -- 14123 FREE #<CONS 0 14124>
 "00000000000000000011011100101101", -- 14124 FREE #<CONS 0 14125>
 "00000000000000000011011100101110", -- 14125 FREE #<CONS 0 14126>
 "00000000000000000011011100101111", -- 14126 FREE #<CONS 0 14127>
 "00000000000000000011011100110000", -- 14127 FREE #<CONS 0 14128>
 "00000000000000000011011100110001", -- 14128 FREE #<CONS 0 14129>
 "00000000000000000011011100110010", -- 14129 FREE #<CONS 0 14130>
 "00000000000000000011011100110011", -- 14130 FREE #<CONS 0 14131>
 "00000000000000000011011100110100", -- 14131 FREE #<CONS 0 14132>
 "00000000000000000011011100110101", -- 14132 FREE #<CONS 0 14133>
 "00000000000000000011011100110110", -- 14133 FREE #<CONS 0 14134>
 "00000000000000000011011100110111", -- 14134 FREE #<CONS 0 14135>
 "00000000000000000011011100111000", -- 14135 FREE #<CONS 0 14136>
 "00000000000000000011011100111001", -- 14136 FREE #<CONS 0 14137>
 "00000000000000000011011100111010", -- 14137 FREE #<CONS 0 14138>
 "00000000000000000011011100111011", -- 14138 FREE #<CONS 0 14139>
 "00000000000000000011011100111100", -- 14139 FREE #<CONS 0 14140>
 "00000000000000000011011100111101", -- 14140 FREE #<CONS 0 14141>
 "00000000000000000011011100111110", -- 14141 FREE #<CONS 0 14142>
 "00000000000000000011011100111111", -- 14142 FREE #<CONS 0 14143>
 "00000000000000000011011101000000", -- 14143 FREE #<CONS 0 14144>
 "00000000000000000011011101000001", -- 14144 FREE #<CONS 0 14145>
 "00000000000000000011011101000010", -- 14145 FREE #<CONS 0 14146>
 "00000000000000000011011101000011", -- 14146 FREE #<CONS 0 14147>
 "00000000000000000011011101000100", -- 14147 FREE #<CONS 0 14148>
 "00000000000000000011011101000101", -- 14148 FREE #<CONS 0 14149>
 "00000000000000000011011101000110", -- 14149 FREE #<CONS 0 14150>
 "00000000000000000011011101000111", -- 14150 FREE #<CONS 0 14151>
 "00000000000000000011011101001000", -- 14151 FREE #<CONS 0 14152>
 "00000000000000000011011101001001", -- 14152 FREE #<CONS 0 14153>
 "00000000000000000011011101001010", -- 14153 FREE #<CONS 0 14154>
 "00000000000000000011011101001011", -- 14154 FREE #<CONS 0 14155>
 "00000000000000000011011101001100", -- 14155 FREE #<CONS 0 14156>
 "00000000000000000011011101001101", -- 14156 FREE #<CONS 0 14157>
 "00000000000000000011011101001110", -- 14157 FREE #<CONS 0 14158>
 "00000000000000000011011101001111", -- 14158 FREE #<CONS 0 14159>
 "00000000000000000011011101010000", -- 14159 FREE #<CONS 0 14160>
 "00000000000000000011011101010001", -- 14160 FREE #<CONS 0 14161>
 "00000000000000000011011101010010", -- 14161 FREE #<CONS 0 14162>
 "00000000000000000011011101010011", -- 14162 FREE #<CONS 0 14163>
 "00000000000000000011011101010100", -- 14163 FREE #<CONS 0 14164>
 "00000000000000000011011101010101", -- 14164 FREE #<CONS 0 14165>
 "00000000000000000011011101010110", -- 14165 FREE #<CONS 0 14166>
 "00000000000000000011011101010111", -- 14166 FREE #<CONS 0 14167>
 "00000000000000000011011101011000", -- 14167 FREE #<CONS 0 14168>
 "00000000000000000011011101011001", -- 14168 FREE #<CONS 0 14169>
 "00000000000000000011011101011010", -- 14169 FREE #<CONS 0 14170>
 "00000000000000000011011101011011", -- 14170 FREE #<CONS 0 14171>
 "00000000000000000011011101011100", -- 14171 FREE #<CONS 0 14172>
 "00000000000000000011011101011101", -- 14172 FREE #<CONS 0 14173>
 "00000000000000000011011101011110", -- 14173 FREE #<CONS 0 14174>
 "00000000000000000011011101011111", -- 14174 FREE #<CONS 0 14175>
 "00000000000000000011011101100000", -- 14175 FREE #<CONS 0 14176>
 "00000000000000000011011101100001", -- 14176 FREE #<CONS 0 14177>
 "00000000000000000011011101100010", -- 14177 FREE #<CONS 0 14178>
 "00000000000000000011011101100011", -- 14178 FREE #<CONS 0 14179>
 "00000000000000000011011101100100", -- 14179 FREE #<CONS 0 14180>
 "00000000000000000011011101100101", -- 14180 FREE #<CONS 0 14181>
 "00000000000000000011011101100110", -- 14181 FREE #<CONS 0 14182>
 "00000000000000000011011101100111", -- 14182 FREE #<CONS 0 14183>
 "00000000000000000011011101101000", -- 14183 FREE #<CONS 0 14184>
 "00000000000000000011011101101001", -- 14184 FREE #<CONS 0 14185>
 "00000000000000000011011101101010", -- 14185 FREE #<CONS 0 14186>
 "00000000000000000011011101101011", -- 14186 FREE #<CONS 0 14187>
 "00000000000000000011011101101100", -- 14187 FREE #<CONS 0 14188>
 "00000000000000000011011101101101", -- 14188 FREE #<CONS 0 14189>
 "00000000000000000011011101101110", -- 14189 FREE #<CONS 0 14190>
 "00000000000000000011011101101111", -- 14190 FREE #<CONS 0 14191>
 "00000000000000000011011101110000", -- 14191 FREE #<CONS 0 14192>
 "00000000000000000011011101110001", -- 14192 FREE #<CONS 0 14193>
 "00000000000000000011011101110010", -- 14193 FREE #<CONS 0 14194>
 "00000000000000000011011101110011", -- 14194 FREE #<CONS 0 14195>
 "00000000000000000011011101110100", -- 14195 FREE #<CONS 0 14196>
 "00000000000000000011011101110101", -- 14196 FREE #<CONS 0 14197>
 "00000000000000000011011101110110", -- 14197 FREE #<CONS 0 14198>
 "00000000000000000011011101110111", -- 14198 FREE #<CONS 0 14199>
 "00000000000000000011011101111000", -- 14199 FREE #<CONS 0 14200>
 "00000000000000000011011101111001", -- 14200 FREE #<CONS 0 14201>
 "00000000000000000011011101111010", -- 14201 FREE #<CONS 0 14202>
 "00000000000000000011011101111011", -- 14202 FREE #<CONS 0 14203>
 "00000000000000000011011101111100", -- 14203 FREE #<CONS 0 14204>
 "00000000000000000011011101111101", -- 14204 FREE #<CONS 0 14205>
 "00000000000000000011011101111110", -- 14205 FREE #<CONS 0 14206>
 "00000000000000000011011101111111", -- 14206 FREE #<CONS 0 14207>
 "00000000000000000011011110000000", -- 14207 FREE #<CONS 0 14208>
 "00000000000000000011011110000001", -- 14208 FREE #<CONS 0 14209>
 "00000000000000000011011110000010", -- 14209 FREE #<CONS 0 14210>
 "00000000000000000011011110000011", -- 14210 FREE #<CONS 0 14211>
 "00000000000000000011011110000100", -- 14211 FREE #<CONS 0 14212>
 "00000000000000000011011110000101", -- 14212 FREE #<CONS 0 14213>
 "00000000000000000011011110000110", -- 14213 FREE #<CONS 0 14214>
 "00000000000000000011011110000111", -- 14214 FREE #<CONS 0 14215>
 "00000000000000000011011110001000", -- 14215 FREE #<CONS 0 14216>
 "00000000000000000011011110001001", -- 14216 FREE #<CONS 0 14217>
 "00000000000000000011011110001010", -- 14217 FREE #<CONS 0 14218>
 "00000000000000000011011110001011", -- 14218 FREE #<CONS 0 14219>
 "00000000000000000011011110001100", -- 14219 FREE #<CONS 0 14220>
 "00000000000000000011011110001101", -- 14220 FREE #<CONS 0 14221>
 "00000000000000000011011110001110", -- 14221 FREE #<CONS 0 14222>
 "00000000000000000011011110001111", -- 14222 FREE #<CONS 0 14223>
 "00000000000000000011011110010000", -- 14223 FREE #<CONS 0 14224>
 "00000000000000000011011110010001", -- 14224 FREE #<CONS 0 14225>
 "00000000000000000011011110010010", -- 14225 FREE #<CONS 0 14226>
 "00000000000000000011011110010011", -- 14226 FREE #<CONS 0 14227>
 "00000000000000000011011110010100", -- 14227 FREE #<CONS 0 14228>
 "00000000000000000011011110010101", -- 14228 FREE #<CONS 0 14229>
 "00000000000000000011011110010110", -- 14229 FREE #<CONS 0 14230>
 "00000000000000000011011110010111", -- 14230 FREE #<CONS 0 14231>
 "00000000000000000011011110011000", -- 14231 FREE #<CONS 0 14232>
 "00000000000000000011011110011001", -- 14232 FREE #<CONS 0 14233>
 "00000000000000000011011110011010", -- 14233 FREE #<CONS 0 14234>
 "00000000000000000011011110011011", -- 14234 FREE #<CONS 0 14235>
 "00000000000000000011011110011100", -- 14235 FREE #<CONS 0 14236>
 "00000000000000000011011110011101", -- 14236 FREE #<CONS 0 14237>
 "00000000000000000011011110011110", -- 14237 FREE #<CONS 0 14238>
 "00000000000000000011011110011111", -- 14238 FREE #<CONS 0 14239>
 "00000000000000000011011110100000", -- 14239 FREE #<CONS 0 14240>
 "00000000000000000011011110100001", -- 14240 FREE #<CONS 0 14241>
 "00000000000000000011011110100010", -- 14241 FREE #<CONS 0 14242>
 "00000000000000000011011110100011", -- 14242 FREE #<CONS 0 14243>
 "00000000000000000011011110100100", -- 14243 FREE #<CONS 0 14244>
 "00000000000000000011011110100101", -- 14244 FREE #<CONS 0 14245>
 "00000000000000000011011110100110", -- 14245 FREE #<CONS 0 14246>
 "00000000000000000011011110100111", -- 14246 FREE #<CONS 0 14247>
 "00000000000000000011011110101000", -- 14247 FREE #<CONS 0 14248>
 "00000000000000000011011110101001", -- 14248 FREE #<CONS 0 14249>
 "00000000000000000011011110101010", -- 14249 FREE #<CONS 0 14250>
 "00000000000000000011011110101011", -- 14250 FREE #<CONS 0 14251>
 "00000000000000000011011110101100", -- 14251 FREE #<CONS 0 14252>
 "00000000000000000011011110101101", -- 14252 FREE #<CONS 0 14253>
 "00000000000000000011011110101110", -- 14253 FREE #<CONS 0 14254>
 "00000000000000000011011110101111", -- 14254 FREE #<CONS 0 14255>
 "00000000000000000011011110110000", -- 14255 FREE #<CONS 0 14256>
 "00000000000000000011011110110001", -- 14256 FREE #<CONS 0 14257>
 "00000000000000000011011110110010", -- 14257 FREE #<CONS 0 14258>
 "00000000000000000011011110110011", -- 14258 FREE #<CONS 0 14259>
 "00000000000000000011011110110100", -- 14259 FREE #<CONS 0 14260>
 "00000000000000000011011110110101", -- 14260 FREE #<CONS 0 14261>
 "00000000000000000011011110110110", -- 14261 FREE #<CONS 0 14262>
 "00000000000000000011011110110111", -- 14262 FREE #<CONS 0 14263>
 "00000000000000000011011110111000", -- 14263 FREE #<CONS 0 14264>
 "00000000000000000011011110111001", -- 14264 FREE #<CONS 0 14265>
 "00000000000000000011011110111010", -- 14265 FREE #<CONS 0 14266>
 "00000000000000000011011110111011", -- 14266 FREE #<CONS 0 14267>
 "00000000000000000011011110111100", -- 14267 FREE #<CONS 0 14268>
 "00000000000000000011011110111101", -- 14268 FREE #<CONS 0 14269>
 "00000000000000000011011110111110", -- 14269 FREE #<CONS 0 14270>
 "00000000000000000011011110111111", -- 14270 FREE #<CONS 0 14271>
 "00000000000000000011011111000000", -- 14271 FREE #<CONS 0 14272>
 "00000000000000000011011111000001", -- 14272 FREE #<CONS 0 14273>
 "00000000000000000011011111000010", -- 14273 FREE #<CONS 0 14274>
 "00000000000000000011011111000011", -- 14274 FREE #<CONS 0 14275>
 "00000000000000000011011111000100", -- 14275 FREE #<CONS 0 14276>
 "00000000000000000011011111000101", -- 14276 FREE #<CONS 0 14277>
 "00000000000000000011011111000110", -- 14277 FREE #<CONS 0 14278>
 "00000000000000000011011111000111", -- 14278 FREE #<CONS 0 14279>
 "00000000000000000011011111001000", -- 14279 FREE #<CONS 0 14280>
 "00000000000000000011011111001001", -- 14280 FREE #<CONS 0 14281>
 "00000000000000000011011111001010", -- 14281 FREE #<CONS 0 14282>
 "00000000000000000011011111001011", -- 14282 FREE #<CONS 0 14283>
 "00000000000000000011011111001100", -- 14283 FREE #<CONS 0 14284>
 "00000000000000000011011111001101", -- 14284 FREE #<CONS 0 14285>
 "00000000000000000011011111001110", -- 14285 FREE #<CONS 0 14286>
 "00000000000000000011011111001111", -- 14286 FREE #<CONS 0 14287>
 "00000000000000000011011111010000", -- 14287 FREE #<CONS 0 14288>
 "00000000000000000011011111010001", -- 14288 FREE #<CONS 0 14289>
 "00000000000000000011011111010010", -- 14289 FREE #<CONS 0 14290>
 "00000000000000000011011111010011", -- 14290 FREE #<CONS 0 14291>
 "00000000000000000011011111010100", -- 14291 FREE #<CONS 0 14292>
 "00000000000000000011011111010101", -- 14292 FREE #<CONS 0 14293>
 "00000000000000000011011111010110", -- 14293 FREE #<CONS 0 14294>
 "00000000000000000011011111010111", -- 14294 FREE #<CONS 0 14295>
 "00000000000000000011011111011000", -- 14295 FREE #<CONS 0 14296>
 "00000000000000000011011111011001", -- 14296 FREE #<CONS 0 14297>
 "00000000000000000011011111011010", -- 14297 FREE #<CONS 0 14298>
 "00000000000000000011011111011011", -- 14298 FREE #<CONS 0 14299>
 "00000000000000000011011111011100", -- 14299 FREE #<CONS 0 14300>
 "00000000000000000011011111011101", -- 14300 FREE #<CONS 0 14301>
 "00000000000000000011011111011110", -- 14301 FREE #<CONS 0 14302>
 "00000000000000000011011111011111", -- 14302 FREE #<CONS 0 14303>
 "00000000000000000011011111100000", -- 14303 FREE #<CONS 0 14304>
 "00000000000000000011011111100001", -- 14304 FREE #<CONS 0 14305>
 "00000000000000000011011111100010", -- 14305 FREE #<CONS 0 14306>
 "00000000000000000011011111100011", -- 14306 FREE #<CONS 0 14307>
 "00000000000000000011011111100100", -- 14307 FREE #<CONS 0 14308>
 "00000000000000000011011111100101", -- 14308 FREE #<CONS 0 14309>
 "00000000000000000011011111100110", -- 14309 FREE #<CONS 0 14310>
 "00000000000000000011011111100111", -- 14310 FREE #<CONS 0 14311>
 "00000000000000000011011111101000", -- 14311 FREE #<CONS 0 14312>
 "00000000000000000011011111101001", -- 14312 FREE #<CONS 0 14313>
 "00000000000000000011011111101010", -- 14313 FREE #<CONS 0 14314>
 "00000000000000000011011111101011", -- 14314 FREE #<CONS 0 14315>
 "00000000000000000011011111101100", -- 14315 FREE #<CONS 0 14316>
 "00000000000000000011011111101101", -- 14316 FREE #<CONS 0 14317>
 "00000000000000000011011111101110", -- 14317 FREE #<CONS 0 14318>
 "00000000000000000011011111101111", -- 14318 FREE #<CONS 0 14319>
 "00000000000000000011011111110000", -- 14319 FREE #<CONS 0 14320>
 "00000000000000000011011111110001", -- 14320 FREE #<CONS 0 14321>
 "00000000000000000011011111110010", -- 14321 FREE #<CONS 0 14322>
 "00000000000000000011011111110011", -- 14322 FREE #<CONS 0 14323>
 "00000000000000000011011111110100", -- 14323 FREE #<CONS 0 14324>
 "00000000000000000011011111110101", -- 14324 FREE #<CONS 0 14325>
 "00000000000000000011011111110110", -- 14325 FREE #<CONS 0 14326>
 "00000000000000000011011111110111", -- 14326 FREE #<CONS 0 14327>
 "00000000000000000011011111111000", -- 14327 FREE #<CONS 0 14328>
 "00000000000000000011011111111001", -- 14328 FREE #<CONS 0 14329>
 "00000000000000000011011111111010", -- 14329 FREE #<CONS 0 14330>
 "00000000000000000011011111111011", -- 14330 FREE #<CONS 0 14331>
 "00000000000000000011011111111100", -- 14331 FREE #<CONS 0 14332>
 "00000000000000000011011111111101", -- 14332 FREE #<CONS 0 14333>
 "00000000000000000011011111111110", -- 14333 FREE #<CONS 0 14334>
 "00000000000000000011011111111111", -- 14334 FREE #<CONS 0 14335>
 "00000000000000000011100000000000", -- 14335 FREE #<CONS 0 14336>
 "00000000000000000011100000000001", -- 14336 FREE #<CONS 0 14337>
 "00000000000000000011100000000010", -- 14337 FREE #<CONS 0 14338>
 "00000000000000000011100000000011", -- 14338 FREE #<CONS 0 14339>
 "00000000000000000011100000000100", -- 14339 FREE #<CONS 0 14340>
 "00000000000000000011100000000101", -- 14340 FREE #<CONS 0 14341>
 "00000000000000000011100000000110", -- 14341 FREE #<CONS 0 14342>
 "00000000000000000011100000000111", -- 14342 FREE #<CONS 0 14343>
 "00000000000000000011100000001000", -- 14343 FREE #<CONS 0 14344>
 "00000000000000000011100000001001", -- 14344 FREE #<CONS 0 14345>
 "00000000000000000011100000001010", -- 14345 FREE #<CONS 0 14346>
 "00000000000000000011100000001011", -- 14346 FREE #<CONS 0 14347>
 "00000000000000000011100000001100", -- 14347 FREE #<CONS 0 14348>
 "00000000000000000011100000001101", -- 14348 FREE #<CONS 0 14349>
 "00000000000000000011100000001110", -- 14349 FREE #<CONS 0 14350>
 "00000000000000000011100000001111", -- 14350 FREE #<CONS 0 14351>
 "00000000000000000011100000010000", -- 14351 FREE #<CONS 0 14352>
 "00000000000000000011100000010001", -- 14352 FREE #<CONS 0 14353>
 "00000000000000000011100000010010", -- 14353 FREE #<CONS 0 14354>
 "00000000000000000011100000010011", -- 14354 FREE #<CONS 0 14355>
 "00000000000000000011100000010100", -- 14355 FREE #<CONS 0 14356>
 "00000000000000000011100000010101", -- 14356 FREE #<CONS 0 14357>
 "00000000000000000011100000010110", -- 14357 FREE #<CONS 0 14358>
 "00000000000000000011100000010111", -- 14358 FREE #<CONS 0 14359>
 "00000000000000000011100000011000", -- 14359 FREE #<CONS 0 14360>
 "00000000000000000011100000011001", -- 14360 FREE #<CONS 0 14361>
 "00000000000000000011100000011010", -- 14361 FREE #<CONS 0 14362>
 "00000000000000000011100000011011", -- 14362 FREE #<CONS 0 14363>
 "00000000000000000011100000011100", -- 14363 FREE #<CONS 0 14364>
 "00000000000000000011100000011101", -- 14364 FREE #<CONS 0 14365>
 "00000000000000000011100000011110", -- 14365 FREE #<CONS 0 14366>
 "00000000000000000011100000011111", -- 14366 FREE #<CONS 0 14367>
 "00000000000000000011100000100000", -- 14367 FREE #<CONS 0 14368>
 "00000000000000000011100000100001", -- 14368 FREE #<CONS 0 14369>
 "00000000000000000011100000100010", -- 14369 FREE #<CONS 0 14370>
 "00000000000000000011100000100011", -- 14370 FREE #<CONS 0 14371>
 "00000000000000000011100000100100", -- 14371 FREE #<CONS 0 14372>
 "00000000000000000011100000100101", -- 14372 FREE #<CONS 0 14373>
 "00000000000000000011100000100110", -- 14373 FREE #<CONS 0 14374>
 "00000000000000000011100000100111", -- 14374 FREE #<CONS 0 14375>
 "00000000000000000011100000101000", -- 14375 FREE #<CONS 0 14376>
 "00000000000000000011100000101001", -- 14376 FREE #<CONS 0 14377>
 "00000000000000000011100000101010", -- 14377 FREE #<CONS 0 14378>
 "00000000000000000011100000101011", -- 14378 FREE #<CONS 0 14379>
 "00000000000000000011100000101100", -- 14379 FREE #<CONS 0 14380>
 "00000000000000000011100000101101", -- 14380 FREE #<CONS 0 14381>
 "00000000000000000011100000101110", -- 14381 FREE #<CONS 0 14382>
 "00000000000000000011100000101111", -- 14382 FREE #<CONS 0 14383>
 "00000000000000000011100000110000", -- 14383 FREE #<CONS 0 14384>
 "00000000000000000011100000110001", -- 14384 FREE #<CONS 0 14385>
 "00000000000000000011100000110010", -- 14385 FREE #<CONS 0 14386>
 "00000000000000000011100000110011", -- 14386 FREE #<CONS 0 14387>
 "00000000000000000011100000110100", -- 14387 FREE #<CONS 0 14388>
 "00000000000000000011100000110101", -- 14388 FREE #<CONS 0 14389>
 "00000000000000000011100000110110", -- 14389 FREE #<CONS 0 14390>
 "00000000000000000011100000110111", -- 14390 FREE #<CONS 0 14391>
 "00000000000000000011100000111000", -- 14391 FREE #<CONS 0 14392>
 "00000000000000000011100000111001", -- 14392 FREE #<CONS 0 14393>
 "00000000000000000011100000111010", -- 14393 FREE #<CONS 0 14394>
 "00000000000000000011100000111011", -- 14394 FREE #<CONS 0 14395>
 "00000000000000000011100000111100", -- 14395 FREE #<CONS 0 14396>
 "00000000000000000011100000111101", -- 14396 FREE #<CONS 0 14397>
 "00000000000000000011100000111110", -- 14397 FREE #<CONS 0 14398>
 "00000000000000000011100000111111", -- 14398 FREE #<CONS 0 14399>
 "00000000000000000011100001000000", -- 14399 FREE #<CONS 0 14400>
 "00000000000000000011100001000001", -- 14400 FREE #<CONS 0 14401>
 "00000000000000000011100001000010", -- 14401 FREE #<CONS 0 14402>
 "00000000000000000011100001000011", -- 14402 FREE #<CONS 0 14403>
 "00000000000000000011100001000100", -- 14403 FREE #<CONS 0 14404>
 "00000000000000000011100001000101", -- 14404 FREE #<CONS 0 14405>
 "00000000000000000011100001000110", -- 14405 FREE #<CONS 0 14406>
 "00000000000000000011100001000111", -- 14406 FREE #<CONS 0 14407>
 "00000000000000000011100001001000", -- 14407 FREE #<CONS 0 14408>
 "00000000000000000011100001001001", -- 14408 FREE #<CONS 0 14409>
 "00000000000000000011100001001010", -- 14409 FREE #<CONS 0 14410>
 "00000000000000000011100001001011", -- 14410 FREE #<CONS 0 14411>
 "00000000000000000011100001001100", -- 14411 FREE #<CONS 0 14412>
 "00000000000000000011100001001101", -- 14412 FREE #<CONS 0 14413>
 "00000000000000000011100001001110", -- 14413 FREE #<CONS 0 14414>
 "00000000000000000011100001001111", -- 14414 FREE #<CONS 0 14415>
 "00000000000000000011100001010000", -- 14415 FREE #<CONS 0 14416>
 "00000000000000000011100001010001", -- 14416 FREE #<CONS 0 14417>
 "00000000000000000011100001010010", -- 14417 FREE #<CONS 0 14418>
 "00000000000000000011100001010011", -- 14418 FREE #<CONS 0 14419>
 "00000000000000000011100001010100", -- 14419 FREE #<CONS 0 14420>
 "00000000000000000011100001010101", -- 14420 FREE #<CONS 0 14421>
 "00000000000000000011100001010110", -- 14421 FREE #<CONS 0 14422>
 "00000000000000000011100001010111", -- 14422 FREE #<CONS 0 14423>
 "00000000000000000011100001011000", -- 14423 FREE #<CONS 0 14424>
 "00000000000000000011100001011001", -- 14424 FREE #<CONS 0 14425>
 "00000000000000000011100001011010", -- 14425 FREE #<CONS 0 14426>
 "00000000000000000011100001011011", -- 14426 FREE #<CONS 0 14427>
 "00000000000000000011100001011100", -- 14427 FREE #<CONS 0 14428>
 "00000000000000000011100001011101", -- 14428 FREE #<CONS 0 14429>
 "00000000000000000011100001011110", -- 14429 FREE #<CONS 0 14430>
 "00000000000000000011100001011111", -- 14430 FREE #<CONS 0 14431>
 "00000000000000000011100001100000", -- 14431 FREE #<CONS 0 14432>
 "00000000000000000011100001100001", -- 14432 FREE #<CONS 0 14433>
 "00000000000000000011100001100010", -- 14433 FREE #<CONS 0 14434>
 "00000000000000000011100001100011", -- 14434 FREE #<CONS 0 14435>
 "00000000000000000011100001100100", -- 14435 FREE #<CONS 0 14436>
 "00000000000000000011100001100101", -- 14436 FREE #<CONS 0 14437>
 "00000000000000000011100001100110", -- 14437 FREE #<CONS 0 14438>
 "00000000000000000011100001100111", -- 14438 FREE #<CONS 0 14439>
 "00000000000000000011100001101000", -- 14439 FREE #<CONS 0 14440>
 "00000000000000000011100001101001", -- 14440 FREE #<CONS 0 14441>
 "00000000000000000011100001101010", -- 14441 FREE #<CONS 0 14442>
 "00000000000000000011100001101011", -- 14442 FREE #<CONS 0 14443>
 "00000000000000000011100001101100", -- 14443 FREE #<CONS 0 14444>
 "00000000000000000011100001101101", -- 14444 FREE #<CONS 0 14445>
 "00000000000000000011100001101110", -- 14445 FREE #<CONS 0 14446>
 "00000000000000000011100001101111", -- 14446 FREE #<CONS 0 14447>
 "00000000000000000011100001110000", -- 14447 FREE #<CONS 0 14448>
 "00000000000000000011100001110001", -- 14448 FREE #<CONS 0 14449>
 "00000000000000000011100001110010", -- 14449 FREE #<CONS 0 14450>
 "00000000000000000011100001110011", -- 14450 FREE #<CONS 0 14451>
 "00000000000000000011100001110100", -- 14451 FREE #<CONS 0 14452>
 "00000000000000000011100001110101", -- 14452 FREE #<CONS 0 14453>
 "00000000000000000011100001110110", -- 14453 FREE #<CONS 0 14454>
 "00000000000000000011100001110111", -- 14454 FREE #<CONS 0 14455>
 "00000000000000000011100001111000", -- 14455 FREE #<CONS 0 14456>
 "00000000000000000011100001111001", -- 14456 FREE #<CONS 0 14457>
 "00000000000000000011100001111010", -- 14457 FREE #<CONS 0 14458>
 "00000000000000000011100001111011", -- 14458 FREE #<CONS 0 14459>
 "00000000000000000011100001111100", -- 14459 FREE #<CONS 0 14460>
 "00000000000000000011100001111101", -- 14460 FREE #<CONS 0 14461>
 "00000000000000000011100001111110", -- 14461 FREE #<CONS 0 14462>
 "00000000000000000011100001111111", -- 14462 FREE #<CONS 0 14463>
 "00000000000000000011100010000000", -- 14463 FREE #<CONS 0 14464>
 "00000000000000000011100010000001", -- 14464 FREE #<CONS 0 14465>
 "00000000000000000011100010000010", -- 14465 FREE #<CONS 0 14466>
 "00000000000000000011100010000011", -- 14466 FREE #<CONS 0 14467>
 "00000000000000000011100010000100", -- 14467 FREE #<CONS 0 14468>
 "00000000000000000011100010000101", -- 14468 FREE #<CONS 0 14469>
 "00000000000000000011100010000110", -- 14469 FREE #<CONS 0 14470>
 "00000000000000000011100010000111", -- 14470 FREE #<CONS 0 14471>
 "00000000000000000011100010001000", -- 14471 FREE #<CONS 0 14472>
 "00000000000000000011100010001001", -- 14472 FREE #<CONS 0 14473>
 "00000000000000000011100010001010", -- 14473 FREE #<CONS 0 14474>
 "00000000000000000011100010001011", -- 14474 FREE #<CONS 0 14475>
 "00000000000000000011100010001100", -- 14475 FREE #<CONS 0 14476>
 "00000000000000000011100010001101", -- 14476 FREE #<CONS 0 14477>
 "00000000000000000011100010001110", -- 14477 FREE #<CONS 0 14478>
 "00000000000000000011100010001111", -- 14478 FREE #<CONS 0 14479>
 "00000000000000000011100010010000", -- 14479 FREE #<CONS 0 14480>
 "00000000000000000011100010010001", -- 14480 FREE #<CONS 0 14481>
 "00000000000000000011100010010010", -- 14481 FREE #<CONS 0 14482>
 "00000000000000000011100010010011", -- 14482 FREE #<CONS 0 14483>
 "00000000000000000011100010010100", -- 14483 FREE #<CONS 0 14484>
 "00000000000000000011100010010101", -- 14484 FREE #<CONS 0 14485>
 "00000000000000000011100010010110", -- 14485 FREE #<CONS 0 14486>
 "00000000000000000011100010010111", -- 14486 FREE #<CONS 0 14487>
 "00000000000000000011100010011000", -- 14487 FREE #<CONS 0 14488>
 "00000000000000000011100010011001", -- 14488 FREE #<CONS 0 14489>
 "00000000000000000011100010011010", -- 14489 FREE #<CONS 0 14490>
 "00000000000000000011100010011011", -- 14490 FREE #<CONS 0 14491>
 "00000000000000000011100010011100", -- 14491 FREE #<CONS 0 14492>
 "00000000000000000011100010011101", -- 14492 FREE #<CONS 0 14493>
 "00000000000000000011100010011110", -- 14493 FREE #<CONS 0 14494>
 "00000000000000000011100010011111", -- 14494 FREE #<CONS 0 14495>
 "00000000000000000011100010100000", -- 14495 FREE #<CONS 0 14496>
 "00000000000000000011100010100001", -- 14496 FREE #<CONS 0 14497>
 "00000000000000000011100010100010", -- 14497 FREE #<CONS 0 14498>
 "00000000000000000011100010100011", -- 14498 FREE #<CONS 0 14499>
 "00000000000000000011100010100100", -- 14499 FREE #<CONS 0 14500>
 "00000000000000000011100010100101", -- 14500 FREE #<CONS 0 14501>
 "00000000000000000011100010100110", -- 14501 FREE #<CONS 0 14502>
 "00000000000000000011100010100111", -- 14502 FREE #<CONS 0 14503>
 "00000000000000000011100010101000", -- 14503 FREE #<CONS 0 14504>
 "00000000000000000011100010101001", -- 14504 FREE #<CONS 0 14505>
 "00000000000000000011100010101010", -- 14505 FREE #<CONS 0 14506>
 "00000000000000000011100010101011", -- 14506 FREE #<CONS 0 14507>
 "00000000000000000011100010101100", -- 14507 FREE #<CONS 0 14508>
 "00000000000000000011100010101101", -- 14508 FREE #<CONS 0 14509>
 "00000000000000000011100010101110", -- 14509 FREE #<CONS 0 14510>
 "00000000000000000011100010101111", -- 14510 FREE #<CONS 0 14511>
 "00000000000000000011100010110000", -- 14511 FREE #<CONS 0 14512>
 "00000000000000000011100010110001", -- 14512 FREE #<CONS 0 14513>
 "00000000000000000011100010110010", -- 14513 FREE #<CONS 0 14514>
 "00000000000000000011100010110011", -- 14514 FREE #<CONS 0 14515>
 "00000000000000000011100010110100", -- 14515 FREE #<CONS 0 14516>
 "00000000000000000011100010110101", -- 14516 FREE #<CONS 0 14517>
 "00000000000000000011100010110110", -- 14517 FREE #<CONS 0 14518>
 "00000000000000000011100010110111", -- 14518 FREE #<CONS 0 14519>
 "00000000000000000011100010111000", -- 14519 FREE #<CONS 0 14520>
 "00000000000000000011100010111001", -- 14520 FREE #<CONS 0 14521>
 "00000000000000000011100010111010", -- 14521 FREE #<CONS 0 14522>
 "00000000000000000011100010111011", -- 14522 FREE #<CONS 0 14523>
 "00000000000000000011100010111100", -- 14523 FREE #<CONS 0 14524>
 "00000000000000000011100010111101", -- 14524 FREE #<CONS 0 14525>
 "00000000000000000011100010111110", -- 14525 FREE #<CONS 0 14526>
 "00000000000000000011100010111111", -- 14526 FREE #<CONS 0 14527>
 "00000000000000000011100011000000", -- 14527 FREE #<CONS 0 14528>
 "00000000000000000011100011000001", -- 14528 FREE #<CONS 0 14529>
 "00000000000000000011100011000010", -- 14529 FREE #<CONS 0 14530>
 "00000000000000000011100011000011", -- 14530 FREE #<CONS 0 14531>
 "00000000000000000011100011000100", -- 14531 FREE #<CONS 0 14532>
 "00000000000000000011100011000101", -- 14532 FREE #<CONS 0 14533>
 "00000000000000000011100011000110", -- 14533 FREE #<CONS 0 14534>
 "00000000000000000011100011000111", -- 14534 FREE #<CONS 0 14535>
 "00000000000000000011100011001000", -- 14535 FREE #<CONS 0 14536>
 "00000000000000000011100011001001", -- 14536 FREE #<CONS 0 14537>
 "00000000000000000011100011001010", -- 14537 FREE #<CONS 0 14538>
 "00000000000000000011100011001011", -- 14538 FREE #<CONS 0 14539>
 "00000000000000000011100011001100", -- 14539 FREE #<CONS 0 14540>
 "00000000000000000011100011001101", -- 14540 FREE #<CONS 0 14541>
 "00000000000000000011100011001110", -- 14541 FREE #<CONS 0 14542>
 "00000000000000000011100011001111", -- 14542 FREE #<CONS 0 14543>
 "00000000000000000011100011010000", -- 14543 FREE #<CONS 0 14544>
 "00000000000000000011100011010001", -- 14544 FREE #<CONS 0 14545>
 "00000000000000000011100011010010", -- 14545 FREE #<CONS 0 14546>
 "00000000000000000011100011010011", -- 14546 FREE #<CONS 0 14547>
 "00000000000000000011100011010100", -- 14547 FREE #<CONS 0 14548>
 "00000000000000000011100011010101", -- 14548 FREE #<CONS 0 14549>
 "00000000000000000011100011010110", -- 14549 FREE #<CONS 0 14550>
 "00000000000000000011100011010111", -- 14550 FREE #<CONS 0 14551>
 "00000000000000000011100011011000", -- 14551 FREE #<CONS 0 14552>
 "00000000000000000011100011011001", -- 14552 FREE #<CONS 0 14553>
 "00000000000000000011100011011010", -- 14553 FREE #<CONS 0 14554>
 "00000000000000000011100011011011", -- 14554 FREE #<CONS 0 14555>
 "00000000000000000011100011011100", -- 14555 FREE #<CONS 0 14556>
 "00000000000000000011100011011101", -- 14556 FREE #<CONS 0 14557>
 "00000000000000000011100011011110", -- 14557 FREE #<CONS 0 14558>
 "00000000000000000011100011011111", -- 14558 FREE #<CONS 0 14559>
 "00000000000000000011100011100000", -- 14559 FREE #<CONS 0 14560>
 "00000000000000000011100011100001", -- 14560 FREE #<CONS 0 14561>
 "00000000000000000011100011100010", -- 14561 FREE #<CONS 0 14562>
 "00000000000000000011100011100011", -- 14562 FREE #<CONS 0 14563>
 "00000000000000000011100011100100", -- 14563 FREE #<CONS 0 14564>
 "00000000000000000011100011100101", -- 14564 FREE #<CONS 0 14565>
 "00000000000000000011100011100110", -- 14565 FREE #<CONS 0 14566>
 "00000000000000000011100011100111", -- 14566 FREE #<CONS 0 14567>
 "00000000000000000011100011101000", -- 14567 FREE #<CONS 0 14568>
 "00000000000000000011100011101001", -- 14568 FREE #<CONS 0 14569>
 "00000000000000000011100011101010", -- 14569 FREE #<CONS 0 14570>
 "00000000000000000011100011101011", -- 14570 FREE #<CONS 0 14571>
 "00000000000000000011100011101100", -- 14571 FREE #<CONS 0 14572>
 "00000000000000000011100011101101", -- 14572 FREE #<CONS 0 14573>
 "00000000000000000011100011101110", -- 14573 FREE #<CONS 0 14574>
 "00000000000000000011100011101111", -- 14574 FREE #<CONS 0 14575>
 "00000000000000000011100011110000", -- 14575 FREE #<CONS 0 14576>
 "00000000000000000011100011110001", -- 14576 FREE #<CONS 0 14577>
 "00000000000000000011100011110010", -- 14577 FREE #<CONS 0 14578>
 "00000000000000000011100011110011", -- 14578 FREE #<CONS 0 14579>
 "00000000000000000011100011110100", -- 14579 FREE #<CONS 0 14580>
 "00000000000000000011100011110101", -- 14580 FREE #<CONS 0 14581>
 "00000000000000000011100011110110", -- 14581 FREE #<CONS 0 14582>
 "00000000000000000011100011110111", -- 14582 FREE #<CONS 0 14583>
 "00000000000000000011100011111000", -- 14583 FREE #<CONS 0 14584>
 "00000000000000000011100011111001", -- 14584 FREE #<CONS 0 14585>
 "00000000000000000011100011111010", -- 14585 FREE #<CONS 0 14586>
 "00000000000000000011100011111011", -- 14586 FREE #<CONS 0 14587>
 "00000000000000000011100011111100", -- 14587 FREE #<CONS 0 14588>
 "00000000000000000011100011111101", -- 14588 FREE #<CONS 0 14589>
 "00000000000000000011100011111110", -- 14589 FREE #<CONS 0 14590>
 "00000000000000000011100011111111", -- 14590 FREE #<CONS 0 14591>
 "00000000000000000011100100000000", -- 14591 FREE #<CONS 0 14592>
 "00000000000000000011100100000001", -- 14592 FREE #<CONS 0 14593>
 "00000000000000000011100100000010", -- 14593 FREE #<CONS 0 14594>
 "00000000000000000011100100000011", -- 14594 FREE #<CONS 0 14595>
 "00000000000000000011100100000100", -- 14595 FREE #<CONS 0 14596>
 "00000000000000000011100100000101", -- 14596 FREE #<CONS 0 14597>
 "00000000000000000011100100000110", -- 14597 FREE #<CONS 0 14598>
 "00000000000000000011100100000111", -- 14598 FREE #<CONS 0 14599>
 "00000000000000000011100100001000", -- 14599 FREE #<CONS 0 14600>
 "00000000000000000011100100001001", -- 14600 FREE #<CONS 0 14601>
 "00000000000000000011100100001010", -- 14601 FREE #<CONS 0 14602>
 "00000000000000000011100100001011", -- 14602 FREE #<CONS 0 14603>
 "00000000000000000011100100001100", -- 14603 FREE #<CONS 0 14604>
 "00000000000000000011100100001101", -- 14604 FREE #<CONS 0 14605>
 "00000000000000000011100100001110", -- 14605 FREE #<CONS 0 14606>
 "00000000000000000011100100001111", -- 14606 FREE #<CONS 0 14607>
 "00000000000000000011100100010000", -- 14607 FREE #<CONS 0 14608>
 "00000000000000000011100100010001", -- 14608 FREE #<CONS 0 14609>
 "00000000000000000011100100010010", -- 14609 FREE #<CONS 0 14610>
 "00000000000000000011100100010011", -- 14610 FREE #<CONS 0 14611>
 "00000000000000000011100100010100", -- 14611 FREE #<CONS 0 14612>
 "00000000000000000011100100010101", -- 14612 FREE #<CONS 0 14613>
 "00000000000000000011100100010110", -- 14613 FREE #<CONS 0 14614>
 "00000000000000000011100100010111", -- 14614 FREE #<CONS 0 14615>
 "00000000000000000011100100011000", -- 14615 FREE #<CONS 0 14616>
 "00000000000000000011100100011001", -- 14616 FREE #<CONS 0 14617>
 "00000000000000000011100100011010", -- 14617 FREE #<CONS 0 14618>
 "00000000000000000011100100011011", -- 14618 FREE #<CONS 0 14619>
 "00000000000000000011100100011100", -- 14619 FREE #<CONS 0 14620>
 "00000000000000000011100100011101", -- 14620 FREE #<CONS 0 14621>
 "00000000000000000011100100011110", -- 14621 FREE #<CONS 0 14622>
 "00000000000000000011100100011111", -- 14622 FREE #<CONS 0 14623>
 "00000000000000000011100100100000", -- 14623 FREE #<CONS 0 14624>
 "00000000000000000011100100100001", -- 14624 FREE #<CONS 0 14625>
 "00000000000000000011100100100010", -- 14625 FREE #<CONS 0 14626>
 "00000000000000000011100100100011", -- 14626 FREE #<CONS 0 14627>
 "00000000000000000011100100100100", -- 14627 FREE #<CONS 0 14628>
 "00000000000000000011100100100101", -- 14628 FREE #<CONS 0 14629>
 "00000000000000000011100100100110", -- 14629 FREE #<CONS 0 14630>
 "00000000000000000011100100100111", -- 14630 FREE #<CONS 0 14631>
 "00000000000000000011100100101000", -- 14631 FREE #<CONS 0 14632>
 "00000000000000000011100100101001", -- 14632 FREE #<CONS 0 14633>
 "00000000000000000011100100101010", -- 14633 FREE #<CONS 0 14634>
 "00000000000000000011100100101011", -- 14634 FREE #<CONS 0 14635>
 "00000000000000000011100100101100", -- 14635 FREE #<CONS 0 14636>
 "00000000000000000011100100101101", -- 14636 FREE #<CONS 0 14637>
 "00000000000000000011100100101110", -- 14637 FREE #<CONS 0 14638>
 "00000000000000000011100100101111", -- 14638 FREE #<CONS 0 14639>
 "00000000000000000011100100110000", -- 14639 FREE #<CONS 0 14640>
 "00000000000000000011100100110001", -- 14640 FREE #<CONS 0 14641>
 "00000000000000000011100100110010", -- 14641 FREE #<CONS 0 14642>
 "00000000000000000011100100110011", -- 14642 FREE #<CONS 0 14643>
 "00000000000000000011100100110100", -- 14643 FREE #<CONS 0 14644>
 "00000000000000000011100100110101", -- 14644 FREE #<CONS 0 14645>
 "00000000000000000011100100110110", -- 14645 FREE #<CONS 0 14646>
 "00000000000000000011100100110111", -- 14646 FREE #<CONS 0 14647>
 "00000000000000000011100100111000", -- 14647 FREE #<CONS 0 14648>
 "00000000000000000011100100111001", -- 14648 FREE #<CONS 0 14649>
 "00000000000000000011100100111010", -- 14649 FREE #<CONS 0 14650>
 "00000000000000000011100100111011", -- 14650 FREE #<CONS 0 14651>
 "00000000000000000011100100111100", -- 14651 FREE #<CONS 0 14652>
 "00000000000000000011100100111101", -- 14652 FREE #<CONS 0 14653>
 "00000000000000000011100100111110", -- 14653 FREE #<CONS 0 14654>
 "00000000000000000011100100111111", -- 14654 FREE #<CONS 0 14655>
 "00000000000000000011100101000000", -- 14655 FREE #<CONS 0 14656>
 "00000000000000000011100101000001", -- 14656 FREE #<CONS 0 14657>
 "00000000000000000011100101000010", -- 14657 FREE #<CONS 0 14658>
 "00000000000000000011100101000011", -- 14658 FREE #<CONS 0 14659>
 "00000000000000000011100101000100", -- 14659 FREE #<CONS 0 14660>
 "00000000000000000011100101000101", -- 14660 FREE #<CONS 0 14661>
 "00000000000000000011100101000110", -- 14661 FREE #<CONS 0 14662>
 "00000000000000000011100101000111", -- 14662 FREE #<CONS 0 14663>
 "00000000000000000011100101001000", -- 14663 FREE #<CONS 0 14664>
 "00000000000000000011100101001001", -- 14664 FREE #<CONS 0 14665>
 "00000000000000000011100101001010", -- 14665 FREE #<CONS 0 14666>
 "00000000000000000011100101001011", -- 14666 FREE #<CONS 0 14667>
 "00000000000000000011100101001100", -- 14667 FREE #<CONS 0 14668>
 "00000000000000000011100101001101", -- 14668 FREE #<CONS 0 14669>
 "00000000000000000011100101001110", -- 14669 FREE #<CONS 0 14670>
 "00000000000000000011100101001111", -- 14670 FREE #<CONS 0 14671>
 "00000000000000000011100101010000", -- 14671 FREE #<CONS 0 14672>
 "00000000000000000011100101010001", -- 14672 FREE #<CONS 0 14673>
 "00000000000000000011100101010010", -- 14673 FREE #<CONS 0 14674>
 "00000000000000000011100101010011", -- 14674 FREE #<CONS 0 14675>
 "00000000000000000011100101010100", -- 14675 FREE #<CONS 0 14676>
 "00000000000000000011100101010101", -- 14676 FREE #<CONS 0 14677>
 "00000000000000000011100101010110", -- 14677 FREE #<CONS 0 14678>
 "00000000000000000011100101010111", -- 14678 FREE #<CONS 0 14679>
 "00000000000000000011100101011000", -- 14679 FREE #<CONS 0 14680>
 "00000000000000000011100101011001", -- 14680 FREE #<CONS 0 14681>
 "00000000000000000011100101011010", -- 14681 FREE #<CONS 0 14682>
 "00000000000000000011100101011011", -- 14682 FREE #<CONS 0 14683>
 "00000000000000000011100101011100", -- 14683 FREE #<CONS 0 14684>
 "00000000000000000011100101011101", -- 14684 FREE #<CONS 0 14685>
 "00000000000000000011100101011110", -- 14685 FREE #<CONS 0 14686>
 "00000000000000000011100101011111", -- 14686 FREE #<CONS 0 14687>
 "00000000000000000011100101100000", -- 14687 FREE #<CONS 0 14688>
 "00000000000000000011100101100001", -- 14688 FREE #<CONS 0 14689>
 "00000000000000000011100101100010", -- 14689 FREE #<CONS 0 14690>
 "00000000000000000011100101100011", -- 14690 FREE #<CONS 0 14691>
 "00000000000000000011100101100100", -- 14691 FREE #<CONS 0 14692>
 "00000000000000000011100101100101", -- 14692 FREE #<CONS 0 14693>
 "00000000000000000011100101100110", -- 14693 FREE #<CONS 0 14694>
 "00000000000000000011100101100111", -- 14694 FREE #<CONS 0 14695>
 "00000000000000000011100101101000", -- 14695 FREE #<CONS 0 14696>
 "00000000000000000011100101101001", -- 14696 FREE #<CONS 0 14697>
 "00000000000000000011100101101010", -- 14697 FREE #<CONS 0 14698>
 "00000000000000000011100101101011", -- 14698 FREE #<CONS 0 14699>
 "00000000000000000011100101101100", -- 14699 FREE #<CONS 0 14700>
 "00000000000000000011100101101101", -- 14700 FREE #<CONS 0 14701>
 "00000000000000000011100101101110", -- 14701 FREE #<CONS 0 14702>
 "00000000000000000011100101101111", -- 14702 FREE #<CONS 0 14703>
 "00000000000000000011100101110000", -- 14703 FREE #<CONS 0 14704>
 "00000000000000000011100101110001", -- 14704 FREE #<CONS 0 14705>
 "00000000000000000011100101110010", -- 14705 FREE #<CONS 0 14706>
 "00000000000000000011100101110011", -- 14706 FREE #<CONS 0 14707>
 "00000000000000000011100101110100", -- 14707 FREE #<CONS 0 14708>
 "00000000000000000011100101110101", -- 14708 FREE #<CONS 0 14709>
 "00000000000000000011100101110110", -- 14709 FREE #<CONS 0 14710>
 "00000000000000000011100101110111", -- 14710 FREE #<CONS 0 14711>
 "00000000000000000011100101111000", -- 14711 FREE #<CONS 0 14712>
 "00000000000000000011100101111001", -- 14712 FREE #<CONS 0 14713>
 "00000000000000000011100101111010", -- 14713 FREE #<CONS 0 14714>
 "00000000000000000011100101111011", -- 14714 FREE #<CONS 0 14715>
 "00000000000000000011100101111100", -- 14715 FREE #<CONS 0 14716>
 "00000000000000000011100101111101", -- 14716 FREE #<CONS 0 14717>
 "00000000000000000011100101111110", -- 14717 FREE #<CONS 0 14718>
 "00000000000000000011100101111111", -- 14718 FREE #<CONS 0 14719>
 "00000000000000000011100110000000", -- 14719 FREE #<CONS 0 14720>
 "00000000000000000011100110000001", -- 14720 FREE #<CONS 0 14721>
 "00000000000000000011100110000010", -- 14721 FREE #<CONS 0 14722>
 "00000000000000000011100110000011", -- 14722 FREE #<CONS 0 14723>
 "00000000000000000011100110000100", -- 14723 FREE #<CONS 0 14724>
 "00000000000000000011100110000101", -- 14724 FREE #<CONS 0 14725>
 "00000000000000000011100110000110", -- 14725 FREE #<CONS 0 14726>
 "00000000000000000011100110000111", -- 14726 FREE #<CONS 0 14727>
 "00000000000000000011100110001000", -- 14727 FREE #<CONS 0 14728>
 "00000000000000000011100110001001", -- 14728 FREE #<CONS 0 14729>
 "00000000000000000011100110001010", -- 14729 FREE #<CONS 0 14730>
 "00000000000000000011100110001011", -- 14730 FREE #<CONS 0 14731>
 "00000000000000000011100110001100", -- 14731 FREE #<CONS 0 14732>
 "00000000000000000011100110001101", -- 14732 FREE #<CONS 0 14733>
 "00000000000000000011100110001110", -- 14733 FREE #<CONS 0 14734>
 "00000000000000000011100110001111", -- 14734 FREE #<CONS 0 14735>
 "00000000000000000011100110010000", -- 14735 FREE #<CONS 0 14736>
 "00000000000000000011100110010001", -- 14736 FREE #<CONS 0 14737>
 "00000000000000000011100110010010", -- 14737 FREE #<CONS 0 14738>
 "00000000000000000011100110010011", -- 14738 FREE #<CONS 0 14739>
 "00000000000000000011100110010100", -- 14739 FREE #<CONS 0 14740>
 "00000000000000000011100110010101", -- 14740 FREE #<CONS 0 14741>
 "00000000000000000011100110010110", -- 14741 FREE #<CONS 0 14742>
 "00000000000000000011100110010111", -- 14742 FREE #<CONS 0 14743>
 "00000000000000000011100110011000", -- 14743 FREE #<CONS 0 14744>
 "00000000000000000011100110011001", -- 14744 FREE #<CONS 0 14745>
 "00000000000000000011100110011010", -- 14745 FREE #<CONS 0 14746>
 "00000000000000000011100110011011", -- 14746 FREE #<CONS 0 14747>
 "00000000000000000011100110011100", -- 14747 FREE #<CONS 0 14748>
 "00000000000000000011100110011101", -- 14748 FREE #<CONS 0 14749>
 "00000000000000000011100110011110", -- 14749 FREE #<CONS 0 14750>
 "00000000000000000011100110011111", -- 14750 FREE #<CONS 0 14751>
 "00000000000000000011100110100000", -- 14751 FREE #<CONS 0 14752>
 "00000000000000000011100110100001", -- 14752 FREE #<CONS 0 14753>
 "00000000000000000011100110100010", -- 14753 FREE #<CONS 0 14754>
 "00000000000000000011100110100011", -- 14754 FREE #<CONS 0 14755>
 "00000000000000000011100110100100", -- 14755 FREE #<CONS 0 14756>
 "00000000000000000011100110100101", -- 14756 FREE #<CONS 0 14757>
 "00000000000000000011100110100110", -- 14757 FREE #<CONS 0 14758>
 "00000000000000000011100110100111", -- 14758 FREE #<CONS 0 14759>
 "00000000000000000011100110101000", -- 14759 FREE #<CONS 0 14760>
 "00000000000000000011100110101001", -- 14760 FREE #<CONS 0 14761>
 "00000000000000000011100110101010", -- 14761 FREE #<CONS 0 14762>
 "00000000000000000011100110101011", -- 14762 FREE #<CONS 0 14763>
 "00000000000000000011100110101100", -- 14763 FREE #<CONS 0 14764>
 "00000000000000000011100110101101", -- 14764 FREE #<CONS 0 14765>
 "00000000000000000011100110101110", -- 14765 FREE #<CONS 0 14766>
 "00000000000000000011100110101111", -- 14766 FREE #<CONS 0 14767>
 "00000000000000000011100110110000", -- 14767 FREE #<CONS 0 14768>
 "00000000000000000011100110110001", -- 14768 FREE #<CONS 0 14769>
 "00000000000000000011100110110010", -- 14769 FREE #<CONS 0 14770>
 "00000000000000000011100110110011", -- 14770 FREE #<CONS 0 14771>
 "00000000000000000011100110110100", -- 14771 FREE #<CONS 0 14772>
 "00000000000000000011100110110101", -- 14772 FREE #<CONS 0 14773>
 "00000000000000000011100110110110", -- 14773 FREE #<CONS 0 14774>
 "00000000000000000011100110110111", -- 14774 FREE #<CONS 0 14775>
 "00000000000000000011100110111000", -- 14775 FREE #<CONS 0 14776>
 "00000000000000000011100110111001", -- 14776 FREE #<CONS 0 14777>
 "00000000000000000011100110111010", -- 14777 FREE #<CONS 0 14778>
 "00000000000000000011100110111011", -- 14778 FREE #<CONS 0 14779>
 "00000000000000000011100110111100", -- 14779 FREE #<CONS 0 14780>
 "00000000000000000011100110111101", -- 14780 FREE #<CONS 0 14781>
 "00000000000000000011100110111110", -- 14781 FREE #<CONS 0 14782>
 "00000000000000000011100110111111", -- 14782 FREE #<CONS 0 14783>
 "00000000000000000011100111000000", -- 14783 FREE #<CONS 0 14784>
 "00000000000000000011100111000001", -- 14784 FREE #<CONS 0 14785>
 "00000000000000000011100111000010", -- 14785 FREE #<CONS 0 14786>
 "00000000000000000011100111000011", -- 14786 FREE #<CONS 0 14787>
 "00000000000000000011100111000100", -- 14787 FREE #<CONS 0 14788>
 "00000000000000000011100111000101", -- 14788 FREE #<CONS 0 14789>
 "00000000000000000011100111000110", -- 14789 FREE #<CONS 0 14790>
 "00000000000000000011100111000111", -- 14790 FREE #<CONS 0 14791>
 "00000000000000000011100111001000", -- 14791 FREE #<CONS 0 14792>
 "00000000000000000011100111001001", -- 14792 FREE #<CONS 0 14793>
 "00000000000000000011100111001010", -- 14793 FREE #<CONS 0 14794>
 "00000000000000000011100111001011", -- 14794 FREE #<CONS 0 14795>
 "00000000000000000011100111001100", -- 14795 FREE #<CONS 0 14796>
 "00000000000000000011100111001101", -- 14796 FREE #<CONS 0 14797>
 "00000000000000000011100111001110", -- 14797 FREE #<CONS 0 14798>
 "00000000000000000011100111001111", -- 14798 FREE #<CONS 0 14799>
 "00000000000000000011100111010000", -- 14799 FREE #<CONS 0 14800>
 "00000000000000000011100111010001", -- 14800 FREE #<CONS 0 14801>
 "00000000000000000011100111010010", -- 14801 FREE #<CONS 0 14802>
 "00000000000000000011100111010011", -- 14802 FREE #<CONS 0 14803>
 "00000000000000000011100111010100", -- 14803 FREE #<CONS 0 14804>
 "00000000000000000011100111010101", -- 14804 FREE #<CONS 0 14805>
 "00000000000000000011100111010110", -- 14805 FREE #<CONS 0 14806>
 "00000000000000000011100111010111", -- 14806 FREE #<CONS 0 14807>
 "00000000000000000011100111011000", -- 14807 FREE #<CONS 0 14808>
 "00000000000000000011100111011001", -- 14808 FREE #<CONS 0 14809>
 "00000000000000000011100111011010", -- 14809 FREE #<CONS 0 14810>
 "00000000000000000011100111011011", -- 14810 FREE #<CONS 0 14811>
 "00000000000000000011100111011100", -- 14811 FREE #<CONS 0 14812>
 "00000000000000000011100111011101", -- 14812 FREE #<CONS 0 14813>
 "00000000000000000011100111011110", -- 14813 FREE #<CONS 0 14814>
 "00000000000000000011100111011111", -- 14814 FREE #<CONS 0 14815>
 "00000000000000000011100111100000", -- 14815 FREE #<CONS 0 14816>
 "00000000000000000011100111100001", -- 14816 FREE #<CONS 0 14817>
 "00000000000000000011100111100010", -- 14817 FREE #<CONS 0 14818>
 "00000000000000000011100111100011", -- 14818 FREE #<CONS 0 14819>
 "00000000000000000011100111100100", -- 14819 FREE #<CONS 0 14820>
 "00000000000000000011100111100101", -- 14820 FREE #<CONS 0 14821>
 "00000000000000000011100111100110", -- 14821 FREE #<CONS 0 14822>
 "00000000000000000011100111100111", -- 14822 FREE #<CONS 0 14823>
 "00000000000000000011100111101000", -- 14823 FREE #<CONS 0 14824>
 "00000000000000000011100111101001", -- 14824 FREE #<CONS 0 14825>
 "00000000000000000011100111101010", -- 14825 FREE #<CONS 0 14826>
 "00000000000000000011100111101011", -- 14826 FREE #<CONS 0 14827>
 "00000000000000000011100111101100", -- 14827 FREE #<CONS 0 14828>
 "00000000000000000011100111101101", -- 14828 FREE #<CONS 0 14829>
 "00000000000000000011100111101110", -- 14829 FREE #<CONS 0 14830>
 "00000000000000000011100111101111", -- 14830 FREE #<CONS 0 14831>
 "00000000000000000011100111110000", -- 14831 FREE #<CONS 0 14832>
 "00000000000000000011100111110001", -- 14832 FREE #<CONS 0 14833>
 "00000000000000000011100111110010", -- 14833 FREE #<CONS 0 14834>
 "00000000000000000011100111110011", -- 14834 FREE #<CONS 0 14835>
 "00000000000000000011100111110100", -- 14835 FREE #<CONS 0 14836>
 "00000000000000000011100111110101", -- 14836 FREE #<CONS 0 14837>
 "00000000000000000011100111110110", -- 14837 FREE #<CONS 0 14838>
 "00000000000000000011100111110111", -- 14838 FREE #<CONS 0 14839>
 "00000000000000000011100111111000", -- 14839 FREE #<CONS 0 14840>
 "00000000000000000011100111111001", -- 14840 FREE #<CONS 0 14841>
 "00000000000000000011100111111010", -- 14841 FREE #<CONS 0 14842>
 "00000000000000000011100111111011", -- 14842 FREE #<CONS 0 14843>
 "00000000000000000011100111111100", -- 14843 FREE #<CONS 0 14844>
 "00000000000000000011100111111101", -- 14844 FREE #<CONS 0 14845>
 "00000000000000000011100111111110", -- 14845 FREE #<CONS 0 14846>
 "00000000000000000011100111111111", -- 14846 FREE #<CONS 0 14847>
 "00000000000000000011101000000000", -- 14847 FREE #<CONS 0 14848>
 "00000000000000000011101000000001", -- 14848 FREE #<CONS 0 14849>
 "00000000000000000011101000000010", -- 14849 FREE #<CONS 0 14850>
 "00000000000000000011101000000011", -- 14850 FREE #<CONS 0 14851>
 "00000000000000000011101000000100", -- 14851 FREE #<CONS 0 14852>
 "00000000000000000011101000000101", -- 14852 FREE #<CONS 0 14853>
 "00000000000000000011101000000110", -- 14853 FREE #<CONS 0 14854>
 "00000000000000000011101000000111", -- 14854 FREE #<CONS 0 14855>
 "00000000000000000011101000001000", -- 14855 FREE #<CONS 0 14856>
 "00000000000000000011101000001001", -- 14856 FREE #<CONS 0 14857>
 "00000000000000000011101000001010", -- 14857 FREE #<CONS 0 14858>
 "00000000000000000011101000001011", -- 14858 FREE #<CONS 0 14859>
 "00000000000000000011101000001100", -- 14859 FREE #<CONS 0 14860>
 "00000000000000000011101000001101", -- 14860 FREE #<CONS 0 14861>
 "00000000000000000011101000001110", -- 14861 FREE #<CONS 0 14862>
 "00000000000000000011101000001111", -- 14862 FREE #<CONS 0 14863>
 "00000000000000000011101000010000", -- 14863 FREE #<CONS 0 14864>
 "00000000000000000011101000010001", -- 14864 FREE #<CONS 0 14865>
 "00000000000000000011101000010010", -- 14865 FREE #<CONS 0 14866>
 "00000000000000000011101000010011", -- 14866 FREE #<CONS 0 14867>
 "00000000000000000011101000010100", -- 14867 FREE #<CONS 0 14868>
 "00000000000000000011101000010101", -- 14868 FREE #<CONS 0 14869>
 "00000000000000000011101000010110", -- 14869 FREE #<CONS 0 14870>
 "00000000000000000011101000010111", -- 14870 FREE #<CONS 0 14871>
 "00000000000000000011101000011000", -- 14871 FREE #<CONS 0 14872>
 "00000000000000000011101000011001", -- 14872 FREE #<CONS 0 14873>
 "00000000000000000011101000011010", -- 14873 FREE #<CONS 0 14874>
 "00000000000000000011101000011011", -- 14874 FREE #<CONS 0 14875>
 "00000000000000000011101000011100", -- 14875 FREE #<CONS 0 14876>
 "00000000000000000011101000011101", -- 14876 FREE #<CONS 0 14877>
 "00000000000000000011101000011110", -- 14877 FREE #<CONS 0 14878>
 "00000000000000000011101000011111", -- 14878 FREE #<CONS 0 14879>
 "00000000000000000011101000100000", -- 14879 FREE #<CONS 0 14880>
 "00000000000000000011101000100001", -- 14880 FREE #<CONS 0 14881>
 "00000000000000000011101000100010", -- 14881 FREE #<CONS 0 14882>
 "00000000000000000011101000100011", -- 14882 FREE #<CONS 0 14883>
 "00000000000000000011101000100100", -- 14883 FREE #<CONS 0 14884>
 "00000000000000000011101000100101", -- 14884 FREE #<CONS 0 14885>
 "00000000000000000011101000100110", -- 14885 FREE #<CONS 0 14886>
 "00000000000000000011101000100111", -- 14886 FREE #<CONS 0 14887>
 "00000000000000000011101000101000", -- 14887 FREE #<CONS 0 14888>
 "00000000000000000011101000101001", -- 14888 FREE #<CONS 0 14889>
 "00000000000000000011101000101010", -- 14889 FREE #<CONS 0 14890>
 "00000000000000000011101000101011", -- 14890 FREE #<CONS 0 14891>
 "00000000000000000011101000101100", -- 14891 FREE #<CONS 0 14892>
 "00000000000000000011101000101101", -- 14892 FREE #<CONS 0 14893>
 "00000000000000000011101000101110", -- 14893 FREE #<CONS 0 14894>
 "00000000000000000011101000101111", -- 14894 FREE #<CONS 0 14895>
 "00000000000000000011101000110000", -- 14895 FREE #<CONS 0 14896>
 "00000000000000000011101000110001", -- 14896 FREE #<CONS 0 14897>
 "00000000000000000011101000110010", -- 14897 FREE #<CONS 0 14898>
 "00000000000000000011101000110011", -- 14898 FREE #<CONS 0 14899>
 "00000000000000000011101000110100", -- 14899 FREE #<CONS 0 14900>
 "00000000000000000011101000110101", -- 14900 FREE #<CONS 0 14901>
 "00000000000000000011101000110110", -- 14901 FREE #<CONS 0 14902>
 "00000000000000000011101000110111", -- 14902 FREE #<CONS 0 14903>
 "00000000000000000011101000111000", -- 14903 FREE #<CONS 0 14904>
 "00000000000000000011101000111001", -- 14904 FREE #<CONS 0 14905>
 "00000000000000000011101000111010", -- 14905 FREE #<CONS 0 14906>
 "00000000000000000011101000111011", -- 14906 FREE #<CONS 0 14907>
 "00000000000000000011101000111100", -- 14907 FREE #<CONS 0 14908>
 "00000000000000000011101000111101", -- 14908 FREE #<CONS 0 14909>
 "00000000000000000011101000111110", -- 14909 FREE #<CONS 0 14910>
 "00000000000000000011101000111111", -- 14910 FREE #<CONS 0 14911>
 "00000000000000000011101001000000", -- 14911 FREE #<CONS 0 14912>
 "00000000000000000011101001000001", -- 14912 FREE #<CONS 0 14913>
 "00000000000000000011101001000010", -- 14913 FREE #<CONS 0 14914>
 "00000000000000000011101001000011", -- 14914 FREE #<CONS 0 14915>
 "00000000000000000011101001000100", -- 14915 FREE #<CONS 0 14916>
 "00000000000000000011101001000101", -- 14916 FREE #<CONS 0 14917>
 "00000000000000000011101001000110", -- 14917 FREE #<CONS 0 14918>
 "00000000000000000011101001000111", -- 14918 FREE #<CONS 0 14919>
 "00000000000000000011101001001000", -- 14919 FREE #<CONS 0 14920>
 "00000000000000000011101001001001", -- 14920 FREE #<CONS 0 14921>
 "00000000000000000011101001001010", -- 14921 FREE #<CONS 0 14922>
 "00000000000000000011101001001011", -- 14922 FREE #<CONS 0 14923>
 "00000000000000000011101001001100", -- 14923 FREE #<CONS 0 14924>
 "00000000000000000011101001001101", -- 14924 FREE #<CONS 0 14925>
 "00000000000000000011101001001110", -- 14925 FREE #<CONS 0 14926>
 "00000000000000000011101001001111", -- 14926 FREE #<CONS 0 14927>
 "00000000000000000011101001010000", -- 14927 FREE #<CONS 0 14928>
 "00000000000000000011101001010001", -- 14928 FREE #<CONS 0 14929>
 "00000000000000000011101001010010", -- 14929 FREE #<CONS 0 14930>
 "00000000000000000011101001010011", -- 14930 FREE #<CONS 0 14931>
 "00000000000000000011101001010100", -- 14931 FREE #<CONS 0 14932>
 "00000000000000000011101001010101", -- 14932 FREE #<CONS 0 14933>
 "00000000000000000011101001010110", -- 14933 FREE #<CONS 0 14934>
 "00000000000000000011101001010111", -- 14934 FREE #<CONS 0 14935>
 "00000000000000000011101001011000", -- 14935 FREE #<CONS 0 14936>
 "00000000000000000011101001011001", -- 14936 FREE #<CONS 0 14937>
 "00000000000000000011101001011010", -- 14937 FREE #<CONS 0 14938>
 "00000000000000000011101001011011", -- 14938 FREE #<CONS 0 14939>
 "00000000000000000011101001011100", -- 14939 FREE #<CONS 0 14940>
 "00000000000000000011101001011101", -- 14940 FREE #<CONS 0 14941>
 "00000000000000000011101001011110", -- 14941 FREE #<CONS 0 14942>
 "00000000000000000011101001011111", -- 14942 FREE #<CONS 0 14943>
 "00000000000000000011101001100000", -- 14943 FREE #<CONS 0 14944>
 "00000000000000000011101001100001", -- 14944 FREE #<CONS 0 14945>
 "00000000000000000011101001100010", -- 14945 FREE #<CONS 0 14946>
 "00000000000000000011101001100011", -- 14946 FREE #<CONS 0 14947>
 "00000000000000000011101001100100", -- 14947 FREE #<CONS 0 14948>
 "00000000000000000011101001100101", -- 14948 FREE #<CONS 0 14949>
 "00000000000000000011101001100110", -- 14949 FREE #<CONS 0 14950>
 "00000000000000000011101001100111", -- 14950 FREE #<CONS 0 14951>
 "00000000000000000011101001101000", -- 14951 FREE #<CONS 0 14952>
 "00000000000000000011101001101001", -- 14952 FREE #<CONS 0 14953>
 "00000000000000000011101001101010", -- 14953 FREE #<CONS 0 14954>
 "00000000000000000011101001101011", -- 14954 FREE #<CONS 0 14955>
 "00000000000000000011101001101100", -- 14955 FREE #<CONS 0 14956>
 "00000000000000000011101001101101", -- 14956 FREE #<CONS 0 14957>
 "00000000000000000011101001101110", -- 14957 FREE #<CONS 0 14958>
 "00000000000000000011101001101111", -- 14958 FREE #<CONS 0 14959>
 "00000000000000000011101001110000", -- 14959 FREE #<CONS 0 14960>
 "00000000000000000011101001110001", -- 14960 FREE #<CONS 0 14961>
 "00000000000000000011101001110010", -- 14961 FREE #<CONS 0 14962>
 "00000000000000000011101001110011", -- 14962 FREE #<CONS 0 14963>
 "00000000000000000011101001110100", -- 14963 FREE #<CONS 0 14964>
 "00000000000000000011101001110101", -- 14964 FREE #<CONS 0 14965>
 "00000000000000000011101001110110", -- 14965 FREE #<CONS 0 14966>
 "00000000000000000011101001110111", -- 14966 FREE #<CONS 0 14967>
 "00000000000000000011101001111000", -- 14967 FREE #<CONS 0 14968>
 "00000000000000000011101001111001", -- 14968 FREE #<CONS 0 14969>
 "00000000000000000011101001111010", -- 14969 FREE #<CONS 0 14970>
 "00000000000000000011101001111011", -- 14970 FREE #<CONS 0 14971>
 "00000000000000000011101001111100", -- 14971 FREE #<CONS 0 14972>
 "00000000000000000011101001111101", -- 14972 FREE #<CONS 0 14973>
 "00000000000000000011101001111110", -- 14973 FREE #<CONS 0 14974>
 "00000000000000000011101001111111", -- 14974 FREE #<CONS 0 14975>
 "00000000000000000011101010000000", -- 14975 FREE #<CONS 0 14976>
 "00000000000000000011101010000001", -- 14976 FREE #<CONS 0 14977>
 "00000000000000000011101010000010", -- 14977 FREE #<CONS 0 14978>
 "00000000000000000011101010000011", -- 14978 FREE #<CONS 0 14979>
 "00000000000000000011101010000100", -- 14979 FREE #<CONS 0 14980>
 "00000000000000000011101010000101", -- 14980 FREE #<CONS 0 14981>
 "00000000000000000011101010000110", -- 14981 FREE #<CONS 0 14982>
 "00000000000000000011101010000111", -- 14982 FREE #<CONS 0 14983>
 "00000000000000000011101010001000", -- 14983 FREE #<CONS 0 14984>
 "00000000000000000011101010001001", -- 14984 FREE #<CONS 0 14985>
 "00000000000000000011101010001010", -- 14985 FREE #<CONS 0 14986>
 "00000000000000000011101010001011", -- 14986 FREE #<CONS 0 14987>
 "00000000000000000011101010001100", -- 14987 FREE #<CONS 0 14988>
 "00000000000000000011101010001101", -- 14988 FREE #<CONS 0 14989>
 "00000000000000000011101010001110", -- 14989 FREE #<CONS 0 14990>
 "00000000000000000011101010001111", -- 14990 FREE #<CONS 0 14991>
 "00000000000000000011101010010000", -- 14991 FREE #<CONS 0 14992>
 "00000000000000000011101010010001", -- 14992 FREE #<CONS 0 14993>
 "00000000000000000011101010010010", -- 14993 FREE #<CONS 0 14994>
 "00000000000000000011101010010011", -- 14994 FREE #<CONS 0 14995>
 "00000000000000000011101010010100", -- 14995 FREE #<CONS 0 14996>
 "00000000000000000011101010010101", -- 14996 FREE #<CONS 0 14997>
 "00000000000000000011101010010110", -- 14997 FREE #<CONS 0 14998>
 "00000000000000000011101010010111", -- 14998 FREE #<CONS 0 14999>
 "00000000000000000011101010011000", -- 14999 FREE #<CONS 0 15000>
 "00000000000000000011101010011001", -- 15000 FREE #<CONS 0 15001>
 "00000000000000000011101010011010", -- 15001 FREE #<CONS 0 15002>
 "00000000000000000011101010011011", -- 15002 FREE #<CONS 0 15003>
 "00000000000000000011101010011100", -- 15003 FREE #<CONS 0 15004>
 "00000000000000000011101010011101", -- 15004 FREE #<CONS 0 15005>
 "00000000000000000011101010011110", -- 15005 FREE #<CONS 0 15006>
 "00000000000000000011101010011111", -- 15006 FREE #<CONS 0 15007>
 "00000000000000000011101010100000", -- 15007 FREE #<CONS 0 15008>
 "00000000000000000011101010100001", -- 15008 FREE #<CONS 0 15009>
 "00000000000000000011101010100010", -- 15009 FREE #<CONS 0 15010>
 "00000000000000000011101010100011", -- 15010 FREE #<CONS 0 15011>
 "00000000000000000011101010100100", -- 15011 FREE #<CONS 0 15012>
 "00000000000000000011101010100101", -- 15012 FREE #<CONS 0 15013>
 "00000000000000000011101010100110", -- 15013 FREE #<CONS 0 15014>
 "00000000000000000011101010100111", -- 15014 FREE #<CONS 0 15015>
 "00000000000000000011101010101000", -- 15015 FREE #<CONS 0 15016>
 "00000000000000000011101010101001", -- 15016 FREE #<CONS 0 15017>
 "00000000000000000011101010101010", -- 15017 FREE #<CONS 0 15018>
 "00000000000000000011101010101011", -- 15018 FREE #<CONS 0 15019>
 "00000000000000000011101010101100", -- 15019 FREE #<CONS 0 15020>
 "00000000000000000011101010101101", -- 15020 FREE #<CONS 0 15021>
 "00000000000000000011101010101110", -- 15021 FREE #<CONS 0 15022>
 "00000000000000000011101010101111", -- 15022 FREE #<CONS 0 15023>
 "00000000000000000011101010110000", -- 15023 FREE #<CONS 0 15024>
 "00000000000000000011101010110001", -- 15024 FREE #<CONS 0 15025>
 "00000000000000000011101010110010", -- 15025 FREE #<CONS 0 15026>
 "00000000000000000011101010110011", -- 15026 FREE #<CONS 0 15027>
 "00000000000000000011101010110100", -- 15027 FREE #<CONS 0 15028>
 "00000000000000000011101010110101", -- 15028 FREE #<CONS 0 15029>
 "00000000000000000011101010110110", -- 15029 FREE #<CONS 0 15030>
 "00000000000000000011101010110111", -- 15030 FREE #<CONS 0 15031>
 "00000000000000000011101010111000", -- 15031 FREE #<CONS 0 15032>
 "00000000000000000011101010111001", -- 15032 FREE #<CONS 0 15033>
 "00000000000000000011101010111010", -- 15033 FREE #<CONS 0 15034>
 "00000000000000000011101010111011", -- 15034 FREE #<CONS 0 15035>
 "00000000000000000011101010111100", -- 15035 FREE #<CONS 0 15036>
 "00000000000000000011101010111101", -- 15036 FREE #<CONS 0 15037>
 "00000000000000000011101010111110", -- 15037 FREE #<CONS 0 15038>
 "00000000000000000011101010111111", -- 15038 FREE #<CONS 0 15039>
 "00000000000000000011101011000000", -- 15039 FREE #<CONS 0 15040>
 "00000000000000000011101011000001", -- 15040 FREE #<CONS 0 15041>
 "00000000000000000011101011000010", -- 15041 FREE #<CONS 0 15042>
 "00000000000000000011101011000011", -- 15042 FREE #<CONS 0 15043>
 "00000000000000000011101011000100", -- 15043 FREE #<CONS 0 15044>
 "00000000000000000011101011000101", -- 15044 FREE #<CONS 0 15045>
 "00000000000000000011101011000110", -- 15045 FREE #<CONS 0 15046>
 "00000000000000000011101011000111", -- 15046 FREE #<CONS 0 15047>
 "00000000000000000011101011001000", -- 15047 FREE #<CONS 0 15048>
 "00000000000000000011101011001001", -- 15048 FREE #<CONS 0 15049>
 "00000000000000000011101011001010", -- 15049 FREE #<CONS 0 15050>
 "00000000000000000011101011001011", -- 15050 FREE #<CONS 0 15051>
 "00000000000000000011101011001100", -- 15051 FREE #<CONS 0 15052>
 "00000000000000000011101011001101", -- 15052 FREE #<CONS 0 15053>
 "00000000000000000011101011001110", -- 15053 FREE #<CONS 0 15054>
 "00000000000000000011101011001111", -- 15054 FREE #<CONS 0 15055>
 "00000000000000000011101011010000", -- 15055 FREE #<CONS 0 15056>
 "00000000000000000011101011010001", -- 15056 FREE #<CONS 0 15057>
 "00000000000000000011101011010010", -- 15057 FREE #<CONS 0 15058>
 "00000000000000000011101011010011", -- 15058 FREE #<CONS 0 15059>
 "00000000000000000011101011010100", -- 15059 FREE #<CONS 0 15060>
 "00000000000000000011101011010101", -- 15060 FREE #<CONS 0 15061>
 "00000000000000000011101011010110", -- 15061 FREE #<CONS 0 15062>
 "00000000000000000011101011010111", -- 15062 FREE #<CONS 0 15063>
 "00000000000000000011101011011000", -- 15063 FREE #<CONS 0 15064>
 "00000000000000000011101011011001", -- 15064 FREE #<CONS 0 15065>
 "00000000000000000011101011011010", -- 15065 FREE #<CONS 0 15066>
 "00000000000000000011101011011011", -- 15066 FREE #<CONS 0 15067>
 "00000000000000000011101011011100", -- 15067 FREE #<CONS 0 15068>
 "00000000000000000011101011011101", -- 15068 FREE #<CONS 0 15069>
 "00000000000000000011101011011110", -- 15069 FREE #<CONS 0 15070>
 "00000000000000000011101011011111", -- 15070 FREE #<CONS 0 15071>
 "00000000000000000011101011100000", -- 15071 FREE #<CONS 0 15072>
 "00000000000000000011101011100001", -- 15072 FREE #<CONS 0 15073>
 "00000000000000000011101011100010", -- 15073 FREE #<CONS 0 15074>
 "00000000000000000011101011100011", -- 15074 FREE #<CONS 0 15075>
 "00000000000000000011101011100100", -- 15075 FREE #<CONS 0 15076>
 "00000000000000000011101011100101", -- 15076 FREE #<CONS 0 15077>
 "00000000000000000011101011100110", -- 15077 FREE #<CONS 0 15078>
 "00000000000000000011101011100111", -- 15078 FREE #<CONS 0 15079>
 "00000000000000000011101011101000", -- 15079 FREE #<CONS 0 15080>
 "00000000000000000011101011101001", -- 15080 FREE #<CONS 0 15081>
 "00000000000000000011101011101010", -- 15081 FREE #<CONS 0 15082>
 "00000000000000000011101011101011", -- 15082 FREE #<CONS 0 15083>
 "00000000000000000011101011101100", -- 15083 FREE #<CONS 0 15084>
 "00000000000000000011101011101101", -- 15084 FREE #<CONS 0 15085>
 "00000000000000000011101011101110", -- 15085 FREE #<CONS 0 15086>
 "00000000000000000011101011101111", -- 15086 FREE #<CONS 0 15087>
 "00000000000000000011101011110000", -- 15087 FREE #<CONS 0 15088>
 "00000000000000000011101011110001", -- 15088 FREE #<CONS 0 15089>
 "00000000000000000011101011110010", -- 15089 FREE #<CONS 0 15090>
 "00000000000000000011101011110011", -- 15090 FREE #<CONS 0 15091>
 "00000000000000000011101011110100", -- 15091 FREE #<CONS 0 15092>
 "00000000000000000011101011110101", -- 15092 FREE #<CONS 0 15093>
 "00000000000000000011101011110110", -- 15093 FREE #<CONS 0 15094>
 "00000000000000000011101011110111", -- 15094 FREE #<CONS 0 15095>
 "00000000000000000011101011111000", -- 15095 FREE #<CONS 0 15096>
 "00000000000000000011101011111001", -- 15096 FREE #<CONS 0 15097>
 "00000000000000000011101011111010", -- 15097 FREE #<CONS 0 15098>
 "00000000000000000011101011111011", -- 15098 FREE #<CONS 0 15099>
 "00000000000000000011101011111100", -- 15099 FREE #<CONS 0 15100>
 "00000000000000000011101011111101", -- 15100 FREE #<CONS 0 15101>
 "00000000000000000011101011111110", -- 15101 FREE #<CONS 0 15102>
 "00000000000000000011101011111111", -- 15102 FREE #<CONS 0 15103>
 "00000000000000000011101100000000", -- 15103 FREE #<CONS 0 15104>
 "00000000000000000011101100000001", -- 15104 FREE #<CONS 0 15105>
 "00000000000000000011101100000010", -- 15105 FREE #<CONS 0 15106>
 "00000000000000000011101100000011", -- 15106 FREE #<CONS 0 15107>
 "00000000000000000011101100000100", -- 15107 FREE #<CONS 0 15108>
 "00000000000000000011101100000101", -- 15108 FREE #<CONS 0 15109>
 "00000000000000000011101100000110", -- 15109 FREE #<CONS 0 15110>
 "00000000000000000011101100000111", -- 15110 FREE #<CONS 0 15111>
 "00000000000000000011101100001000", -- 15111 FREE #<CONS 0 15112>
 "00000000000000000011101100001001", -- 15112 FREE #<CONS 0 15113>
 "00000000000000000011101100001010", -- 15113 FREE #<CONS 0 15114>
 "00000000000000000011101100001011", -- 15114 FREE #<CONS 0 15115>
 "00000000000000000011101100001100", -- 15115 FREE #<CONS 0 15116>
 "00000000000000000011101100001101", -- 15116 FREE #<CONS 0 15117>
 "00000000000000000011101100001110", -- 15117 FREE #<CONS 0 15118>
 "00000000000000000011101100001111", -- 15118 FREE #<CONS 0 15119>
 "00000000000000000011101100010000", -- 15119 FREE #<CONS 0 15120>
 "00000000000000000011101100010001", -- 15120 FREE #<CONS 0 15121>
 "00000000000000000011101100010010", -- 15121 FREE #<CONS 0 15122>
 "00000000000000000011101100010011", -- 15122 FREE #<CONS 0 15123>
 "00000000000000000011101100010100", -- 15123 FREE #<CONS 0 15124>
 "00000000000000000011101100010101", -- 15124 FREE #<CONS 0 15125>
 "00000000000000000011101100010110", -- 15125 FREE #<CONS 0 15126>
 "00000000000000000011101100010111", -- 15126 FREE #<CONS 0 15127>
 "00000000000000000011101100011000", -- 15127 FREE #<CONS 0 15128>
 "00000000000000000011101100011001", -- 15128 FREE #<CONS 0 15129>
 "00000000000000000011101100011010", -- 15129 FREE #<CONS 0 15130>
 "00000000000000000011101100011011", -- 15130 FREE #<CONS 0 15131>
 "00000000000000000011101100011100", -- 15131 FREE #<CONS 0 15132>
 "00000000000000000011101100011101", -- 15132 FREE #<CONS 0 15133>
 "00000000000000000011101100011110", -- 15133 FREE #<CONS 0 15134>
 "00000000000000000011101100011111", -- 15134 FREE #<CONS 0 15135>
 "00000000000000000011101100100000", -- 15135 FREE #<CONS 0 15136>
 "00000000000000000011101100100001", -- 15136 FREE #<CONS 0 15137>
 "00000000000000000011101100100010", -- 15137 FREE #<CONS 0 15138>
 "00000000000000000011101100100011", -- 15138 FREE #<CONS 0 15139>
 "00000000000000000011101100100100", -- 15139 FREE #<CONS 0 15140>
 "00000000000000000011101100100101", -- 15140 FREE #<CONS 0 15141>
 "00000000000000000011101100100110", -- 15141 FREE #<CONS 0 15142>
 "00000000000000000011101100100111", -- 15142 FREE #<CONS 0 15143>
 "00000000000000000011101100101000", -- 15143 FREE #<CONS 0 15144>
 "00000000000000000011101100101001", -- 15144 FREE #<CONS 0 15145>
 "00000000000000000011101100101010", -- 15145 FREE #<CONS 0 15146>
 "00000000000000000011101100101011", -- 15146 FREE #<CONS 0 15147>
 "00000000000000000011101100101100", -- 15147 FREE #<CONS 0 15148>
 "00000000000000000011101100101101", -- 15148 FREE #<CONS 0 15149>
 "00000000000000000011101100101110", -- 15149 FREE #<CONS 0 15150>
 "00000000000000000011101100101111", -- 15150 FREE #<CONS 0 15151>
 "00000000000000000011101100110000", -- 15151 FREE #<CONS 0 15152>
 "00000000000000000011101100110001", -- 15152 FREE #<CONS 0 15153>
 "00000000000000000011101100110010", -- 15153 FREE #<CONS 0 15154>
 "00000000000000000011101100110011", -- 15154 FREE #<CONS 0 15155>
 "00000000000000000011101100110100", -- 15155 FREE #<CONS 0 15156>
 "00000000000000000011101100110101", -- 15156 FREE #<CONS 0 15157>
 "00000000000000000011101100110110", -- 15157 FREE #<CONS 0 15158>
 "00000000000000000011101100110111", -- 15158 FREE #<CONS 0 15159>
 "00000000000000000011101100111000", -- 15159 FREE #<CONS 0 15160>
 "00000000000000000011101100111001", -- 15160 FREE #<CONS 0 15161>
 "00000000000000000011101100111010", -- 15161 FREE #<CONS 0 15162>
 "00000000000000000011101100111011", -- 15162 FREE #<CONS 0 15163>
 "00000000000000000011101100111100", -- 15163 FREE #<CONS 0 15164>
 "00000000000000000011101100111101", -- 15164 FREE #<CONS 0 15165>
 "00000000000000000011101100111110", -- 15165 FREE #<CONS 0 15166>
 "00000000000000000011101100111111", -- 15166 FREE #<CONS 0 15167>
 "00000000000000000011101101000000", -- 15167 FREE #<CONS 0 15168>
 "00000000000000000011101101000001", -- 15168 FREE #<CONS 0 15169>
 "00000000000000000011101101000010", -- 15169 FREE #<CONS 0 15170>
 "00000000000000000011101101000011", -- 15170 FREE #<CONS 0 15171>
 "00000000000000000011101101000100", -- 15171 FREE #<CONS 0 15172>
 "00000000000000000011101101000101", -- 15172 FREE #<CONS 0 15173>
 "00000000000000000011101101000110", -- 15173 FREE #<CONS 0 15174>
 "00000000000000000011101101000111", -- 15174 FREE #<CONS 0 15175>
 "00000000000000000011101101001000", -- 15175 FREE #<CONS 0 15176>
 "00000000000000000011101101001001", -- 15176 FREE #<CONS 0 15177>
 "00000000000000000011101101001010", -- 15177 FREE #<CONS 0 15178>
 "00000000000000000011101101001011", -- 15178 FREE #<CONS 0 15179>
 "00000000000000000011101101001100", -- 15179 FREE #<CONS 0 15180>
 "00000000000000000011101101001101", -- 15180 FREE #<CONS 0 15181>
 "00000000000000000011101101001110", -- 15181 FREE #<CONS 0 15182>
 "00000000000000000011101101001111", -- 15182 FREE #<CONS 0 15183>
 "00000000000000000011101101010000", -- 15183 FREE #<CONS 0 15184>
 "00000000000000000011101101010001", -- 15184 FREE #<CONS 0 15185>
 "00000000000000000011101101010010", -- 15185 FREE #<CONS 0 15186>
 "00000000000000000011101101010011", -- 15186 FREE #<CONS 0 15187>
 "00000000000000000011101101010100", -- 15187 FREE #<CONS 0 15188>
 "00000000000000000011101101010101", -- 15188 FREE #<CONS 0 15189>
 "00000000000000000011101101010110", -- 15189 FREE #<CONS 0 15190>
 "00000000000000000011101101010111", -- 15190 FREE #<CONS 0 15191>
 "00000000000000000011101101011000", -- 15191 FREE #<CONS 0 15192>
 "00000000000000000011101101011001", -- 15192 FREE #<CONS 0 15193>
 "00000000000000000011101101011010", -- 15193 FREE #<CONS 0 15194>
 "00000000000000000011101101011011", -- 15194 FREE #<CONS 0 15195>
 "00000000000000000011101101011100", -- 15195 FREE #<CONS 0 15196>
 "00000000000000000011101101011101", -- 15196 FREE #<CONS 0 15197>
 "00000000000000000011101101011110", -- 15197 FREE #<CONS 0 15198>
 "00000000000000000011101101011111", -- 15198 FREE #<CONS 0 15199>
 "00000000000000000011101101100000", -- 15199 FREE #<CONS 0 15200>
 "00000000000000000011101101100001", -- 15200 FREE #<CONS 0 15201>
 "00000000000000000011101101100010", -- 15201 FREE #<CONS 0 15202>
 "00000000000000000011101101100011", -- 15202 FREE #<CONS 0 15203>
 "00000000000000000011101101100100", -- 15203 FREE #<CONS 0 15204>
 "00000000000000000011101101100101", -- 15204 FREE #<CONS 0 15205>
 "00000000000000000011101101100110", -- 15205 FREE #<CONS 0 15206>
 "00000000000000000011101101100111", -- 15206 FREE #<CONS 0 15207>
 "00000000000000000011101101101000", -- 15207 FREE #<CONS 0 15208>
 "00000000000000000011101101101001", -- 15208 FREE #<CONS 0 15209>
 "00000000000000000011101101101010", -- 15209 FREE #<CONS 0 15210>
 "00000000000000000011101101101011", -- 15210 FREE #<CONS 0 15211>
 "00000000000000000011101101101100", -- 15211 FREE #<CONS 0 15212>
 "00000000000000000011101101101101", -- 15212 FREE #<CONS 0 15213>
 "00000000000000000011101101101110", -- 15213 FREE #<CONS 0 15214>
 "00000000000000000011101101101111", -- 15214 FREE #<CONS 0 15215>
 "00000000000000000011101101110000", -- 15215 FREE #<CONS 0 15216>
 "00000000000000000011101101110001", -- 15216 FREE #<CONS 0 15217>
 "00000000000000000011101101110010", -- 15217 FREE #<CONS 0 15218>
 "00000000000000000011101101110011", -- 15218 FREE #<CONS 0 15219>
 "00000000000000000011101101110100", -- 15219 FREE #<CONS 0 15220>
 "00000000000000000011101101110101", -- 15220 FREE #<CONS 0 15221>
 "00000000000000000011101101110110", -- 15221 FREE #<CONS 0 15222>
 "00000000000000000011101101110111", -- 15222 FREE #<CONS 0 15223>
 "00000000000000000011101101111000", -- 15223 FREE #<CONS 0 15224>
 "00000000000000000011101101111001", -- 15224 FREE #<CONS 0 15225>
 "00000000000000000011101101111010", -- 15225 FREE #<CONS 0 15226>
 "00000000000000000011101101111011", -- 15226 FREE #<CONS 0 15227>
 "00000000000000000011101101111100", -- 15227 FREE #<CONS 0 15228>
 "00000000000000000011101101111101", -- 15228 FREE #<CONS 0 15229>
 "00000000000000000011101101111110", -- 15229 FREE #<CONS 0 15230>
 "00000000000000000011101101111111", -- 15230 FREE #<CONS 0 15231>
 "00000000000000000011101110000000", -- 15231 FREE #<CONS 0 15232>
 "00000000000000000011101110000001", -- 15232 FREE #<CONS 0 15233>
 "00000000000000000011101110000010", -- 15233 FREE #<CONS 0 15234>
 "00000000000000000011101110000011", -- 15234 FREE #<CONS 0 15235>
 "00000000000000000011101110000100", -- 15235 FREE #<CONS 0 15236>
 "00000000000000000011101110000101", -- 15236 FREE #<CONS 0 15237>
 "00000000000000000011101110000110", -- 15237 FREE #<CONS 0 15238>
 "00000000000000000011101110000111", -- 15238 FREE #<CONS 0 15239>
 "00000000000000000011101110001000", -- 15239 FREE #<CONS 0 15240>
 "00000000000000000011101110001001", -- 15240 FREE #<CONS 0 15241>
 "00000000000000000011101110001010", -- 15241 FREE #<CONS 0 15242>
 "00000000000000000011101110001011", -- 15242 FREE #<CONS 0 15243>
 "00000000000000000011101110001100", -- 15243 FREE #<CONS 0 15244>
 "00000000000000000011101110001101", -- 15244 FREE #<CONS 0 15245>
 "00000000000000000011101110001110", -- 15245 FREE #<CONS 0 15246>
 "00000000000000000011101110001111", -- 15246 FREE #<CONS 0 15247>
 "00000000000000000011101110010000", -- 15247 FREE #<CONS 0 15248>
 "00000000000000000011101110010001", -- 15248 FREE #<CONS 0 15249>
 "00000000000000000011101110010010", -- 15249 FREE #<CONS 0 15250>
 "00000000000000000011101110010011", -- 15250 FREE #<CONS 0 15251>
 "00000000000000000011101110010100", -- 15251 FREE #<CONS 0 15252>
 "00000000000000000011101110010101", -- 15252 FREE #<CONS 0 15253>
 "00000000000000000011101110010110", -- 15253 FREE #<CONS 0 15254>
 "00000000000000000011101110010111", -- 15254 FREE #<CONS 0 15255>
 "00000000000000000011101110011000", -- 15255 FREE #<CONS 0 15256>
 "00000000000000000011101110011001", -- 15256 FREE #<CONS 0 15257>
 "00000000000000000011101110011010", -- 15257 FREE #<CONS 0 15258>
 "00000000000000000011101110011011", -- 15258 FREE #<CONS 0 15259>
 "00000000000000000011101110011100", -- 15259 FREE #<CONS 0 15260>
 "00000000000000000011101110011101", -- 15260 FREE #<CONS 0 15261>
 "00000000000000000011101110011110", -- 15261 FREE #<CONS 0 15262>
 "00000000000000000011101110011111", -- 15262 FREE #<CONS 0 15263>
 "00000000000000000011101110100000", -- 15263 FREE #<CONS 0 15264>
 "00000000000000000011101110100001", -- 15264 FREE #<CONS 0 15265>
 "00000000000000000011101110100010", -- 15265 FREE #<CONS 0 15266>
 "00000000000000000011101110100011", -- 15266 FREE #<CONS 0 15267>
 "00000000000000000011101110100100", -- 15267 FREE #<CONS 0 15268>
 "00000000000000000011101110100101", -- 15268 FREE #<CONS 0 15269>
 "00000000000000000011101110100110", -- 15269 FREE #<CONS 0 15270>
 "00000000000000000011101110100111", -- 15270 FREE #<CONS 0 15271>
 "00000000000000000011101110101000", -- 15271 FREE #<CONS 0 15272>
 "00000000000000000011101110101001", -- 15272 FREE #<CONS 0 15273>
 "00000000000000000011101110101010", -- 15273 FREE #<CONS 0 15274>
 "00000000000000000011101110101011", -- 15274 FREE #<CONS 0 15275>
 "00000000000000000011101110101100", -- 15275 FREE #<CONS 0 15276>
 "00000000000000000011101110101101", -- 15276 FREE #<CONS 0 15277>
 "00000000000000000011101110101110", -- 15277 FREE #<CONS 0 15278>
 "00000000000000000011101110101111", -- 15278 FREE #<CONS 0 15279>
 "00000000000000000011101110110000", -- 15279 FREE #<CONS 0 15280>
 "00000000000000000011101110110001", -- 15280 FREE #<CONS 0 15281>
 "00000000000000000011101110110010", -- 15281 FREE #<CONS 0 15282>
 "00000000000000000011101110110011", -- 15282 FREE #<CONS 0 15283>
 "00000000000000000011101110110100", -- 15283 FREE #<CONS 0 15284>
 "00000000000000000011101110110101", -- 15284 FREE #<CONS 0 15285>
 "00000000000000000011101110110110", -- 15285 FREE #<CONS 0 15286>
 "00000000000000000011101110110111", -- 15286 FREE #<CONS 0 15287>
 "00000000000000000011101110111000", -- 15287 FREE #<CONS 0 15288>
 "00000000000000000011101110111001", -- 15288 FREE #<CONS 0 15289>
 "00000000000000000011101110111010", -- 15289 FREE #<CONS 0 15290>
 "00000000000000000011101110111011", -- 15290 FREE #<CONS 0 15291>
 "00000000000000000011101110111100", -- 15291 FREE #<CONS 0 15292>
 "00000000000000000011101110111101", -- 15292 FREE #<CONS 0 15293>
 "00000000000000000011101110111110", -- 15293 FREE #<CONS 0 15294>
 "00000000000000000011101110111111", -- 15294 FREE #<CONS 0 15295>
 "00000000000000000011101111000000", -- 15295 FREE #<CONS 0 15296>
 "00000000000000000011101111000001", -- 15296 FREE #<CONS 0 15297>
 "00000000000000000011101111000010", -- 15297 FREE #<CONS 0 15298>
 "00000000000000000011101111000011", -- 15298 FREE #<CONS 0 15299>
 "00000000000000000011101111000100", -- 15299 FREE #<CONS 0 15300>
 "00000000000000000011101111000101", -- 15300 FREE #<CONS 0 15301>
 "00000000000000000011101111000110", -- 15301 FREE #<CONS 0 15302>
 "00000000000000000011101111000111", -- 15302 FREE #<CONS 0 15303>
 "00000000000000000011101111001000", -- 15303 FREE #<CONS 0 15304>
 "00000000000000000011101111001001", -- 15304 FREE #<CONS 0 15305>
 "00000000000000000011101111001010", -- 15305 FREE #<CONS 0 15306>
 "00000000000000000011101111001011", -- 15306 FREE #<CONS 0 15307>
 "00000000000000000011101111001100", -- 15307 FREE #<CONS 0 15308>
 "00000000000000000011101111001101", -- 15308 FREE #<CONS 0 15309>
 "00000000000000000011101111001110", -- 15309 FREE #<CONS 0 15310>
 "00000000000000000011101111001111", -- 15310 FREE #<CONS 0 15311>
 "00000000000000000011101111010000", -- 15311 FREE #<CONS 0 15312>
 "00000000000000000011101111010001", -- 15312 FREE #<CONS 0 15313>
 "00000000000000000011101111010010", -- 15313 FREE #<CONS 0 15314>
 "00000000000000000011101111010011", -- 15314 FREE #<CONS 0 15315>
 "00000000000000000011101111010100", -- 15315 FREE #<CONS 0 15316>
 "00000000000000000011101111010101", -- 15316 FREE #<CONS 0 15317>
 "00000000000000000011101111010110", -- 15317 FREE #<CONS 0 15318>
 "00000000000000000011101111010111", -- 15318 FREE #<CONS 0 15319>
 "00000000000000000011101111011000", -- 15319 FREE #<CONS 0 15320>
 "00000000000000000011101111011001", -- 15320 FREE #<CONS 0 15321>
 "00000000000000000011101111011010", -- 15321 FREE #<CONS 0 15322>
 "00000000000000000011101111011011", -- 15322 FREE #<CONS 0 15323>
 "00000000000000000011101111011100", -- 15323 FREE #<CONS 0 15324>
 "00000000000000000011101111011101", -- 15324 FREE #<CONS 0 15325>
 "00000000000000000011101111011110", -- 15325 FREE #<CONS 0 15326>
 "00000000000000000011101111011111", -- 15326 FREE #<CONS 0 15327>
 "00000000000000000011101111100000", -- 15327 FREE #<CONS 0 15328>
 "00000000000000000011101111100001", -- 15328 FREE #<CONS 0 15329>
 "00000000000000000011101111100010", -- 15329 FREE #<CONS 0 15330>
 "00000000000000000011101111100011", -- 15330 FREE #<CONS 0 15331>
 "00000000000000000011101111100100", -- 15331 FREE #<CONS 0 15332>
 "00000000000000000011101111100101", -- 15332 FREE #<CONS 0 15333>
 "00000000000000000011101111100110", -- 15333 FREE #<CONS 0 15334>
 "00000000000000000011101111100111", -- 15334 FREE #<CONS 0 15335>
 "00000000000000000011101111101000", -- 15335 FREE #<CONS 0 15336>
 "00000000000000000011101111101001", -- 15336 FREE #<CONS 0 15337>
 "00000000000000000011101111101010", -- 15337 FREE #<CONS 0 15338>
 "00000000000000000011101111101011", -- 15338 FREE #<CONS 0 15339>
 "00000000000000000011101111101100", -- 15339 FREE #<CONS 0 15340>
 "00000000000000000011101111101101", -- 15340 FREE #<CONS 0 15341>
 "00000000000000000011101111101110", -- 15341 FREE #<CONS 0 15342>
 "00000000000000000011101111101111", -- 15342 FREE #<CONS 0 15343>
 "00000000000000000011101111110000", -- 15343 FREE #<CONS 0 15344>
 "00000000000000000011101111110001", -- 15344 FREE #<CONS 0 15345>
 "00000000000000000011101111110010", -- 15345 FREE #<CONS 0 15346>
 "00000000000000000011101111110011", -- 15346 FREE #<CONS 0 15347>
 "00000000000000000011101111110100", -- 15347 FREE #<CONS 0 15348>
 "00000000000000000011101111110101", -- 15348 FREE #<CONS 0 15349>
 "00000000000000000011101111110110", -- 15349 FREE #<CONS 0 15350>
 "00000000000000000011101111110111", -- 15350 FREE #<CONS 0 15351>
 "00000000000000000011101111111000", -- 15351 FREE #<CONS 0 15352>
 "00000000000000000011101111111001", -- 15352 FREE #<CONS 0 15353>
 "00000000000000000011101111111010", -- 15353 FREE #<CONS 0 15354>
 "00000000000000000011101111111011", -- 15354 FREE #<CONS 0 15355>
 "00000000000000000011101111111100", -- 15355 FREE #<CONS 0 15356>
 "00000000000000000011101111111101", -- 15356 FREE #<CONS 0 15357>
 "00000000000000000011101111111110", -- 15357 FREE #<CONS 0 15358>
 "00000000000000000011101111111111", -- 15358 FREE #<CONS 0 15359>
 "00000000000000000011110000000000", -- 15359 FREE #<CONS 0 15360>
 "00000000000000000011110000000001", -- 15360 FREE #<CONS 0 15361>
 "00000000000000000011110000000010", -- 15361 FREE #<CONS 0 15362>
 "00000000000000000011110000000011", -- 15362 FREE #<CONS 0 15363>
 "00000000000000000011110000000100", -- 15363 FREE #<CONS 0 15364>
 "00000000000000000011110000000101", -- 15364 FREE #<CONS 0 15365>
 "00000000000000000011110000000110", -- 15365 FREE #<CONS 0 15366>
 "00000000000000000011110000000111", -- 15366 FREE #<CONS 0 15367>
 "00000000000000000011110000001000", -- 15367 FREE #<CONS 0 15368>
 "00000000000000000011110000001001", -- 15368 FREE #<CONS 0 15369>
 "00000000000000000011110000001010", -- 15369 FREE #<CONS 0 15370>
 "00000000000000000011110000001011", -- 15370 FREE #<CONS 0 15371>
 "00000000000000000011110000001100", -- 15371 FREE #<CONS 0 15372>
 "00000000000000000011110000001101", -- 15372 FREE #<CONS 0 15373>
 "00000000000000000011110000001110", -- 15373 FREE #<CONS 0 15374>
 "00000000000000000011110000001111", -- 15374 FREE #<CONS 0 15375>
 "00000000000000000011110000010000", -- 15375 FREE #<CONS 0 15376>
 "00000000000000000011110000010001", -- 15376 FREE #<CONS 0 15377>
 "00000000000000000011110000010010", -- 15377 FREE #<CONS 0 15378>
 "00000000000000000011110000010011", -- 15378 FREE #<CONS 0 15379>
 "00000000000000000011110000010100", -- 15379 FREE #<CONS 0 15380>
 "00000000000000000011110000010101", -- 15380 FREE #<CONS 0 15381>
 "00000000000000000011110000010110", -- 15381 FREE #<CONS 0 15382>
 "00000000000000000011110000010111", -- 15382 FREE #<CONS 0 15383>
 "00000000000000000011110000011000", -- 15383 FREE #<CONS 0 15384>
 "00000000000000000011110000011001", -- 15384 FREE #<CONS 0 15385>
 "00000000000000000011110000011010", -- 15385 FREE #<CONS 0 15386>
 "00000000000000000011110000011011", -- 15386 FREE #<CONS 0 15387>
 "00000000000000000011110000011100", -- 15387 FREE #<CONS 0 15388>
 "00000000000000000011110000011101", -- 15388 FREE #<CONS 0 15389>
 "00000000000000000011110000011110", -- 15389 FREE #<CONS 0 15390>
 "00000000000000000011110000011111", -- 15390 FREE #<CONS 0 15391>
 "00000000000000000011110000100000", -- 15391 FREE #<CONS 0 15392>
 "00000000000000000011110000100001", -- 15392 FREE #<CONS 0 15393>
 "00000000000000000011110000100010", -- 15393 FREE #<CONS 0 15394>
 "00000000000000000011110000100011", -- 15394 FREE #<CONS 0 15395>
 "00000000000000000011110000100100", -- 15395 FREE #<CONS 0 15396>
 "00000000000000000011110000100101", -- 15396 FREE #<CONS 0 15397>
 "00000000000000000011110000100110", -- 15397 FREE #<CONS 0 15398>
 "00000000000000000011110000100111", -- 15398 FREE #<CONS 0 15399>
 "00000000000000000011110000101000", -- 15399 FREE #<CONS 0 15400>
 "00000000000000000011110000101001", -- 15400 FREE #<CONS 0 15401>
 "00000000000000000011110000101010", -- 15401 FREE #<CONS 0 15402>
 "00000000000000000011110000101011", -- 15402 FREE #<CONS 0 15403>
 "00000000000000000011110000101100", -- 15403 FREE #<CONS 0 15404>
 "00000000000000000011110000101101", -- 15404 FREE #<CONS 0 15405>
 "00000000000000000011110000101110", -- 15405 FREE #<CONS 0 15406>
 "00000000000000000011110000101111", -- 15406 FREE #<CONS 0 15407>
 "00000000000000000011110000110000", -- 15407 FREE #<CONS 0 15408>
 "00000000000000000011110000110001", -- 15408 FREE #<CONS 0 15409>
 "00000000000000000011110000110010", -- 15409 FREE #<CONS 0 15410>
 "00000000000000000011110000110011", -- 15410 FREE #<CONS 0 15411>
 "00000000000000000011110000110100", -- 15411 FREE #<CONS 0 15412>
 "00000000000000000011110000110101", -- 15412 FREE #<CONS 0 15413>
 "00000000000000000011110000110110", -- 15413 FREE #<CONS 0 15414>
 "00000000000000000011110000110111", -- 15414 FREE #<CONS 0 15415>
 "00000000000000000011110000111000", -- 15415 FREE #<CONS 0 15416>
 "00000000000000000011110000111001", -- 15416 FREE #<CONS 0 15417>
 "00000000000000000011110000111010", -- 15417 FREE #<CONS 0 15418>
 "00000000000000000011110000111011", -- 15418 FREE #<CONS 0 15419>
 "00000000000000000011110000111100", -- 15419 FREE #<CONS 0 15420>
 "00000000000000000011110000111101", -- 15420 FREE #<CONS 0 15421>
 "00000000000000000011110000111110", -- 15421 FREE #<CONS 0 15422>
 "00000000000000000011110000111111", -- 15422 FREE #<CONS 0 15423>
 "00000000000000000011110001000000", -- 15423 FREE #<CONS 0 15424>
 "00000000000000000011110001000001", -- 15424 FREE #<CONS 0 15425>
 "00000000000000000011110001000010", -- 15425 FREE #<CONS 0 15426>
 "00000000000000000011110001000011", -- 15426 FREE #<CONS 0 15427>
 "00000000000000000011110001000100", -- 15427 FREE #<CONS 0 15428>
 "00000000000000000011110001000101", -- 15428 FREE #<CONS 0 15429>
 "00000000000000000011110001000110", -- 15429 FREE #<CONS 0 15430>
 "00000000000000000011110001000111", -- 15430 FREE #<CONS 0 15431>
 "00000000000000000011110001001000", -- 15431 FREE #<CONS 0 15432>
 "00000000000000000011110001001001", -- 15432 FREE #<CONS 0 15433>
 "00000000000000000011110001001010", -- 15433 FREE #<CONS 0 15434>
 "00000000000000000011110001001011", -- 15434 FREE #<CONS 0 15435>
 "00000000000000000011110001001100", -- 15435 FREE #<CONS 0 15436>
 "00000000000000000011110001001101", -- 15436 FREE #<CONS 0 15437>
 "00000000000000000011110001001110", -- 15437 FREE #<CONS 0 15438>
 "00000000000000000011110001001111", -- 15438 FREE #<CONS 0 15439>
 "00000000000000000011110001010000", -- 15439 FREE #<CONS 0 15440>
 "00000000000000000011110001010001", -- 15440 FREE #<CONS 0 15441>
 "00000000000000000011110001010010", -- 15441 FREE #<CONS 0 15442>
 "00000000000000000011110001010011", -- 15442 FREE #<CONS 0 15443>
 "00000000000000000011110001010100", -- 15443 FREE #<CONS 0 15444>
 "00000000000000000011110001010101", -- 15444 FREE #<CONS 0 15445>
 "00000000000000000011110001010110", -- 15445 FREE #<CONS 0 15446>
 "00000000000000000011110001010111", -- 15446 FREE #<CONS 0 15447>
 "00000000000000000011110001011000", -- 15447 FREE #<CONS 0 15448>
 "00000000000000000011110001011001", -- 15448 FREE #<CONS 0 15449>
 "00000000000000000011110001011010", -- 15449 FREE #<CONS 0 15450>
 "00000000000000000011110001011011", -- 15450 FREE #<CONS 0 15451>
 "00000000000000000011110001011100", -- 15451 FREE #<CONS 0 15452>
 "00000000000000000011110001011101", -- 15452 FREE #<CONS 0 15453>
 "00000000000000000011110001011110", -- 15453 FREE #<CONS 0 15454>
 "00000000000000000011110001011111", -- 15454 FREE #<CONS 0 15455>
 "00000000000000000011110001100000", -- 15455 FREE #<CONS 0 15456>
 "00000000000000000011110001100001", -- 15456 FREE #<CONS 0 15457>
 "00000000000000000011110001100010", -- 15457 FREE #<CONS 0 15458>
 "00000000000000000011110001100011", -- 15458 FREE #<CONS 0 15459>
 "00000000000000000011110001100100", -- 15459 FREE #<CONS 0 15460>
 "00000000000000000011110001100101", -- 15460 FREE #<CONS 0 15461>
 "00000000000000000011110001100110", -- 15461 FREE #<CONS 0 15462>
 "00000000000000000011110001100111", -- 15462 FREE #<CONS 0 15463>
 "00000000000000000011110001101000", -- 15463 FREE #<CONS 0 15464>
 "00000000000000000011110001101001", -- 15464 FREE #<CONS 0 15465>
 "00000000000000000011110001101010", -- 15465 FREE #<CONS 0 15466>
 "00000000000000000011110001101011", -- 15466 FREE #<CONS 0 15467>
 "00000000000000000011110001101100", -- 15467 FREE #<CONS 0 15468>
 "00000000000000000011110001101101", -- 15468 FREE #<CONS 0 15469>
 "00000000000000000011110001101110", -- 15469 FREE #<CONS 0 15470>
 "00000000000000000011110001101111", -- 15470 FREE #<CONS 0 15471>
 "00000000000000000011110001110000", -- 15471 FREE #<CONS 0 15472>
 "00000000000000000011110001110001", -- 15472 FREE #<CONS 0 15473>
 "00000000000000000011110001110010", -- 15473 FREE #<CONS 0 15474>
 "00000000000000000011110001110011", -- 15474 FREE #<CONS 0 15475>
 "00000000000000000011110001110100", -- 15475 FREE #<CONS 0 15476>
 "00000000000000000011110001110101", -- 15476 FREE #<CONS 0 15477>
 "00000000000000000011110001110110", -- 15477 FREE #<CONS 0 15478>
 "00000000000000000011110001110111", -- 15478 FREE #<CONS 0 15479>
 "00000000000000000011110001111000", -- 15479 FREE #<CONS 0 15480>
 "00000000000000000011110001111001", -- 15480 FREE #<CONS 0 15481>
 "00000000000000000011110001111010", -- 15481 FREE #<CONS 0 15482>
 "00000000000000000011110001111011", -- 15482 FREE #<CONS 0 15483>
 "00000000000000000011110001111100", -- 15483 FREE #<CONS 0 15484>
 "00000000000000000011110001111101", -- 15484 FREE #<CONS 0 15485>
 "00000000000000000011110001111110", -- 15485 FREE #<CONS 0 15486>
 "00000000000000000011110001111111", -- 15486 FREE #<CONS 0 15487>
 "00000000000000000011110010000000", -- 15487 FREE #<CONS 0 15488>
 "00000000000000000011110010000001", -- 15488 FREE #<CONS 0 15489>
 "00000000000000000011110010000010", -- 15489 FREE #<CONS 0 15490>
 "00000000000000000011110010000011", -- 15490 FREE #<CONS 0 15491>
 "00000000000000000011110010000100", -- 15491 FREE #<CONS 0 15492>
 "00000000000000000011110010000101", -- 15492 FREE #<CONS 0 15493>
 "00000000000000000011110010000110", -- 15493 FREE #<CONS 0 15494>
 "00000000000000000011110010000111", -- 15494 FREE #<CONS 0 15495>
 "00000000000000000011110010001000", -- 15495 FREE #<CONS 0 15496>
 "00000000000000000011110010001001", -- 15496 FREE #<CONS 0 15497>
 "00000000000000000011110010001010", -- 15497 FREE #<CONS 0 15498>
 "00000000000000000011110010001011", -- 15498 FREE #<CONS 0 15499>
 "00000000000000000011110010001100", -- 15499 FREE #<CONS 0 15500>
 "00000000000000000011110010001101", -- 15500 FREE #<CONS 0 15501>
 "00000000000000000011110010001110", -- 15501 FREE #<CONS 0 15502>
 "00000000000000000011110010001111", -- 15502 FREE #<CONS 0 15503>
 "00000000000000000011110010010000", -- 15503 FREE #<CONS 0 15504>
 "00000000000000000011110010010001", -- 15504 FREE #<CONS 0 15505>
 "00000000000000000011110010010010", -- 15505 FREE #<CONS 0 15506>
 "00000000000000000011110010010011", -- 15506 FREE #<CONS 0 15507>
 "00000000000000000011110010010100", -- 15507 FREE #<CONS 0 15508>
 "00000000000000000011110010010101", -- 15508 FREE #<CONS 0 15509>
 "00000000000000000011110010010110", -- 15509 FREE #<CONS 0 15510>
 "00000000000000000011110010010111", -- 15510 FREE #<CONS 0 15511>
 "00000000000000000011110010011000", -- 15511 FREE #<CONS 0 15512>
 "00000000000000000011110010011001", -- 15512 FREE #<CONS 0 15513>
 "00000000000000000011110010011010", -- 15513 FREE #<CONS 0 15514>
 "00000000000000000011110010011011", -- 15514 FREE #<CONS 0 15515>
 "00000000000000000011110010011100", -- 15515 FREE #<CONS 0 15516>
 "00000000000000000011110010011101", -- 15516 FREE #<CONS 0 15517>
 "00000000000000000011110010011110", -- 15517 FREE #<CONS 0 15518>
 "00000000000000000011110010011111", -- 15518 FREE #<CONS 0 15519>
 "00000000000000000011110010100000", -- 15519 FREE #<CONS 0 15520>
 "00000000000000000011110010100001", -- 15520 FREE #<CONS 0 15521>
 "00000000000000000011110010100010", -- 15521 FREE #<CONS 0 15522>
 "00000000000000000011110010100011", -- 15522 FREE #<CONS 0 15523>
 "00000000000000000011110010100100", -- 15523 FREE #<CONS 0 15524>
 "00000000000000000011110010100101", -- 15524 FREE #<CONS 0 15525>
 "00000000000000000011110010100110", -- 15525 FREE #<CONS 0 15526>
 "00000000000000000011110010100111", -- 15526 FREE #<CONS 0 15527>
 "00000000000000000011110010101000", -- 15527 FREE #<CONS 0 15528>
 "00000000000000000011110010101001", -- 15528 FREE #<CONS 0 15529>
 "00000000000000000011110010101010", -- 15529 FREE #<CONS 0 15530>
 "00000000000000000011110010101011", -- 15530 FREE #<CONS 0 15531>
 "00000000000000000011110010101100", -- 15531 FREE #<CONS 0 15532>
 "00000000000000000011110010101101", -- 15532 FREE #<CONS 0 15533>
 "00000000000000000011110010101110", -- 15533 FREE #<CONS 0 15534>
 "00000000000000000011110010101111", -- 15534 FREE #<CONS 0 15535>
 "00000000000000000011110010110000", -- 15535 FREE #<CONS 0 15536>
 "00000000000000000011110010110001", -- 15536 FREE #<CONS 0 15537>
 "00000000000000000011110010110010", -- 15537 FREE #<CONS 0 15538>
 "00000000000000000011110010110011", -- 15538 FREE #<CONS 0 15539>
 "00000000000000000011110010110100", -- 15539 FREE #<CONS 0 15540>
 "00000000000000000011110010110101", -- 15540 FREE #<CONS 0 15541>
 "00000000000000000011110010110110", -- 15541 FREE #<CONS 0 15542>
 "00000000000000000011110010110111", -- 15542 FREE #<CONS 0 15543>
 "00000000000000000011110010111000", -- 15543 FREE #<CONS 0 15544>
 "00000000000000000011110010111001", -- 15544 FREE #<CONS 0 15545>
 "00000000000000000011110010111010", -- 15545 FREE #<CONS 0 15546>
 "00000000000000000011110010111011", -- 15546 FREE #<CONS 0 15547>
 "00000000000000000011110010111100", -- 15547 FREE #<CONS 0 15548>
 "00000000000000000011110010111101", -- 15548 FREE #<CONS 0 15549>
 "00000000000000000011110010111110", -- 15549 FREE #<CONS 0 15550>
 "00000000000000000011110010111111", -- 15550 FREE #<CONS 0 15551>
 "00000000000000000011110011000000", -- 15551 FREE #<CONS 0 15552>
 "00000000000000000011110011000001", -- 15552 FREE #<CONS 0 15553>
 "00000000000000000011110011000010", -- 15553 FREE #<CONS 0 15554>
 "00000000000000000011110011000011", -- 15554 FREE #<CONS 0 15555>
 "00000000000000000011110011000100", -- 15555 FREE #<CONS 0 15556>
 "00000000000000000011110011000101", -- 15556 FREE #<CONS 0 15557>
 "00000000000000000011110011000110", -- 15557 FREE #<CONS 0 15558>
 "00000000000000000011110011000111", -- 15558 FREE #<CONS 0 15559>
 "00000000000000000011110011001000", -- 15559 FREE #<CONS 0 15560>
 "00000000000000000011110011001001", -- 15560 FREE #<CONS 0 15561>
 "00000000000000000011110011001010", -- 15561 FREE #<CONS 0 15562>
 "00000000000000000011110011001011", -- 15562 FREE #<CONS 0 15563>
 "00000000000000000011110011001100", -- 15563 FREE #<CONS 0 15564>
 "00000000000000000011110011001101", -- 15564 FREE #<CONS 0 15565>
 "00000000000000000011110011001110", -- 15565 FREE #<CONS 0 15566>
 "00000000000000000011110011001111", -- 15566 FREE #<CONS 0 15567>
 "00000000000000000011110011010000", -- 15567 FREE #<CONS 0 15568>
 "00000000000000000011110011010001", -- 15568 FREE #<CONS 0 15569>
 "00000000000000000011110011010010", -- 15569 FREE #<CONS 0 15570>
 "00000000000000000011110011010011", -- 15570 FREE #<CONS 0 15571>
 "00000000000000000011110011010100", -- 15571 FREE #<CONS 0 15572>
 "00000000000000000011110011010101", -- 15572 FREE #<CONS 0 15573>
 "00000000000000000011110011010110", -- 15573 FREE #<CONS 0 15574>
 "00000000000000000011110011010111", -- 15574 FREE #<CONS 0 15575>
 "00000000000000000011110011011000", -- 15575 FREE #<CONS 0 15576>
 "00000000000000000011110011011001", -- 15576 FREE #<CONS 0 15577>
 "00000000000000000011110011011010", -- 15577 FREE #<CONS 0 15578>
 "00000000000000000011110011011011", -- 15578 FREE #<CONS 0 15579>
 "00000000000000000011110011011100", -- 15579 FREE #<CONS 0 15580>
 "00000000000000000011110011011101", -- 15580 FREE #<CONS 0 15581>
 "00000000000000000011110011011110", -- 15581 FREE #<CONS 0 15582>
 "00000000000000000011110011011111", -- 15582 FREE #<CONS 0 15583>
 "00000000000000000011110011100000", -- 15583 FREE #<CONS 0 15584>
 "00000000000000000011110011100001", -- 15584 FREE #<CONS 0 15585>
 "00000000000000000011110011100010", -- 15585 FREE #<CONS 0 15586>
 "00000000000000000011110011100011", -- 15586 FREE #<CONS 0 15587>
 "00000000000000000011110011100100", -- 15587 FREE #<CONS 0 15588>
 "00000000000000000011110011100101", -- 15588 FREE #<CONS 0 15589>
 "00000000000000000011110011100110", -- 15589 FREE #<CONS 0 15590>
 "00000000000000000011110011100111", -- 15590 FREE #<CONS 0 15591>
 "00000000000000000011110011101000", -- 15591 FREE #<CONS 0 15592>
 "00000000000000000011110011101001", -- 15592 FREE #<CONS 0 15593>
 "00000000000000000011110011101010", -- 15593 FREE #<CONS 0 15594>
 "00000000000000000011110011101011", -- 15594 FREE #<CONS 0 15595>
 "00000000000000000011110011101100", -- 15595 FREE #<CONS 0 15596>
 "00000000000000000011110011101101", -- 15596 FREE #<CONS 0 15597>
 "00000000000000000011110011101110", -- 15597 FREE #<CONS 0 15598>
 "00000000000000000011110011101111", -- 15598 FREE #<CONS 0 15599>
 "00000000000000000011110011110000", -- 15599 FREE #<CONS 0 15600>
 "00000000000000000011110011110001", -- 15600 FREE #<CONS 0 15601>
 "00000000000000000011110011110010", -- 15601 FREE #<CONS 0 15602>
 "00000000000000000011110011110011", -- 15602 FREE #<CONS 0 15603>
 "00000000000000000011110011110100", -- 15603 FREE #<CONS 0 15604>
 "00000000000000000011110011110101", -- 15604 FREE #<CONS 0 15605>
 "00000000000000000011110011110110", -- 15605 FREE #<CONS 0 15606>
 "00000000000000000011110011110111", -- 15606 FREE #<CONS 0 15607>
 "00000000000000000011110011111000", -- 15607 FREE #<CONS 0 15608>
 "00000000000000000011110011111001", -- 15608 FREE #<CONS 0 15609>
 "00000000000000000011110011111010", -- 15609 FREE #<CONS 0 15610>
 "00000000000000000011110011111011", -- 15610 FREE #<CONS 0 15611>
 "00000000000000000011110011111100", -- 15611 FREE #<CONS 0 15612>
 "00000000000000000011110011111101", -- 15612 FREE #<CONS 0 15613>
 "00000000000000000011110011111110", -- 15613 FREE #<CONS 0 15614>
 "00000000000000000011110011111111", -- 15614 FREE #<CONS 0 15615>
 "00000000000000000011110100000000", -- 15615 FREE #<CONS 0 15616>
 "00000000000000000011110100000001", -- 15616 FREE #<CONS 0 15617>
 "00000000000000000011110100000010", -- 15617 FREE #<CONS 0 15618>
 "00000000000000000011110100000011", -- 15618 FREE #<CONS 0 15619>
 "00000000000000000011110100000100", -- 15619 FREE #<CONS 0 15620>
 "00000000000000000011110100000101", -- 15620 FREE #<CONS 0 15621>
 "00000000000000000011110100000110", -- 15621 FREE #<CONS 0 15622>
 "00000000000000000011110100000111", -- 15622 FREE #<CONS 0 15623>
 "00000000000000000011110100001000", -- 15623 FREE #<CONS 0 15624>
 "00000000000000000011110100001001", -- 15624 FREE #<CONS 0 15625>
 "00000000000000000011110100001010", -- 15625 FREE #<CONS 0 15626>
 "00000000000000000011110100001011", -- 15626 FREE #<CONS 0 15627>
 "00000000000000000011110100001100", -- 15627 FREE #<CONS 0 15628>
 "00000000000000000011110100001101", -- 15628 FREE #<CONS 0 15629>
 "00000000000000000011110100001110", -- 15629 FREE #<CONS 0 15630>
 "00000000000000000011110100001111", -- 15630 FREE #<CONS 0 15631>
 "00000000000000000011110100010000", -- 15631 FREE #<CONS 0 15632>
 "00000000000000000011110100010001", -- 15632 FREE #<CONS 0 15633>
 "00000000000000000011110100010010", -- 15633 FREE #<CONS 0 15634>
 "00000000000000000011110100010011", -- 15634 FREE #<CONS 0 15635>
 "00000000000000000011110100010100", -- 15635 FREE #<CONS 0 15636>
 "00000000000000000011110100010101", -- 15636 FREE #<CONS 0 15637>
 "00000000000000000011110100010110", -- 15637 FREE #<CONS 0 15638>
 "00000000000000000011110100010111", -- 15638 FREE #<CONS 0 15639>
 "00000000000000000011110100011000", -- 15639 FREE #<CONS 0 15640>
 "00000000000000000011110100011001", -- 15640 FREE #<CONS 0 15641>
 "00000000000000000011110100011010", -- 15641 FREE #<CONS 0 15642>
 "00000000000000000011110100011011", -- 15642 FREE #<CONS 0 15643>
 "00000000000000000011110100011100", -- 15643 FREE #<CONS 0 15644>
 "00000000000000000011110100011101", -- 15644 FREE #<CONS 0 15645>
 "00000000000000000011110100011110", -- 15645 FREE #<CONS 0 15646>
 "00000000000000000011110100011111", -- 15646 FREE #<CONS 0 15647>
 "00000000000000000011110100100000", -- 15647 FREE #<CONS 0 15648>
 "00000000000000000011110100100001", -- 15648 FREE #<CONS 0 15649>
 "00000000000000000011110100100010", -- 15649 FREE #<CONS 0 15650>
 "00000000000000000011110100100011", -- 15650 FREE #<CONS 0 15651>
 "00000000000000000011110100100100", -- 15651 FREE #<CONS 0 15652>
 "00000000000000000011110100100101", -- 15652 FREE #<CONS 0 15653>
 "00000000000000000011110100100110", -- 15653 FREE #<CONS 0 15654>
 "00000000000000000011110100100111", -- 15654 FREE #<CONS 0 15655>
 "00000000000000000011110100101000", -- 15655 FREE #<CONS 0 15656>
 "00000000000000000011110100101001", -- 15656 FREE #<CONS 0 15657>
 "00000000000000000011110100101010", -- 15657 FREE #<CONS 0 15658>
 "00000000000000000011110100101011", -- 15658 FREE #<CONS 0 15659>
 "00000000000000000011110100101100", -- 15659 FREE #<CONS 0 15660>
 "00000000000000000011110100101101", -- 15660 FREE #<CONS 0 15661>
 "00000000000000000011110100101110", -- 15661 FREE #<CONS 0 15662>
 "00000000000000000011110100101111", -- 15662 FREE #<CONS 0 15663>
 "00000000000000000011110100110000", -- 15663 FREE #<CONS 0 15664>
 "00000000000000000011110100110001", -- 15664 FREE #<CONS 0 15665>
 "00000000000000000011110100110010", -- 15665 FREE #<CONS 0 15666>
 "00000000000000000011110100110011", -- 15666 FREE #<CONS 0 15667>
 "00000000000000000011110100110100", -- 15667 FREE #<CONS 0 15668>
 "00000000000000000011110100110101", -- 15668 FREE #<CONS 0 15669>
 "00000000000000000011110100110110", -- 15669 FREE #<CONS 0 15670>
 "00000000000000000011110100110111", -- 15670 FREE #<CONS 0 15671>
 "00000000000000000011110100111000", -- 15671 FREE #<CONS 0 15672>
 "00000000000000000011110100111001", -- 15672 FREE #<CONS 0 15673>
 "00000000000000000011110100111010", -- 15673 FREE #<CONS 0 15674>
 "00000000000000000011110100111011", -- 15674 FREE #<CONS 0 15675>
 "00000000000000000011110100111100", -- 15675 FREE #<CONS 0 15676>
 "00000000000000000011110100111101", -- 15676 FREE #<CONS 0 15677>
 "00000000000000000011110100111110", -- 15677 FREE #<CONS 0 15678>
 "00000000000000000011110100111111", -- 15678 FREE #<CONS 0 15679>
 "00000000000000000011110101000000", -- 15679 FREE #<CONS 0 15680>
 "00000000000000000011110101000001", -- 15680 FREE #<CONS 0 15681>
 "00000000000000000011110101000010", -- 15681 FREE #<CONS 0 15682>
 "00000000000000000011110101000011", -- 15682 FREE #<CONS 0 15683>
 "00000000000000000011110101000100", -- 15683 FREE #<CONS 0 15684>
 "00000000000000000011110101000101", -- 15684 FREE #<CONS 0 15685>
 "00000000000000000011110101000110", -- 15685 FREE #<CONS 0 15686>
 "00000000000000000011110101000111", -- 15686 FREE #<CONS 0 15687>
 "00000000000000000011110101001000", -- 15687 FREE #<CONS 0 15688>
 "00000000000000000011110101001001", -- 15688 FREE #<CONS 0 15689>
 "00000000000000000011110101001010", -- 15689 FREE #<CONS 0 15690>
 "00000000000000000011110101001011", -- 15690 FREE #<CONS 0 15691>
 "00000000000000000011110101001100", -- 15691 FREE #<CONS 0 15692>
 "00000000000000000011110101001101", -- 15692 FREE #<CONS 0 15693>
 "00000000000000000011110101001110", -- 15693 FREE #<CONS 0 15694>
 "00000000000000000011110101001111", -- 15694 FREE #<CONS 0 15695>
 "00000000000000000011110101010000", -- 15695 FREE #<CONS 0 15696>
 "00000000000000000011110101010001", -- 15696 FREE #<CONS 0 15697>
 "00000000000000000011110101010010", -- 15697 FREE #<CONS 0 15698>
 "00000000000000000011110101010011", -- 15698 FREE #<CONS 0 15699>
 "00000000000000000011110101010100", -- 15699 FREE #<CONS 0 15700>
 "00000000000000000011110101010101", -- 15700 FREE #<CONS 0 15701>
 "00000000000000000011110101010110", -- 15701 FREE #<CONS 0 15702>
 "00000000000000000011110101010111", -- 15702 FREE #<CONS 0 15703>
 "00000000000000000011110101011000", -- 15703 FREE #<CONS 0 15704>
 "00000000000000000011110101011001", -- 15704 FREE #<CONS 0 15705>
 "00000000000000000011110101011010", -- 15705 FREE #<CONS 0 15706>
 "00000000000000000011110101011011", -- 15706 FREE #<CONS 0 15707>
 "00000000000000000011110101011100", -- 15707 FREE #<CONS 0 15708>
 "00000000000000000011110101011101", -- 15708 FREE #<CONS 0 15709>
 "00000000000000000011110101011110", -- 15709 FREE #<CONS 0 15710>
 "00000000000000000011110101011111", -- 15710 FREE #<CONS 0 15711>
 "00000000000000000011110101100000", -- 15711 FREE #<CONS 0 15712>
 "00000000000000000011110101100001", -- 15712 FREE #<CONS 0 15713>
 "00000000000000000011110101100010", -- 15713 FREE #<CONS 0 15714>
 "00000000000000000011110101100011", -- 15714 FREE #<CONS 0 15715>
 "00000000000000000011110101100100", -- 15715 FREE #<CONS 0 15716>
 "00000000000000000011110101100101", -- 15716 FREE #<CONS 0 15717>
 "00000000000000000011110101100110", -- 15717 FREE #<CONS 0 15718>
 "00000000000000000011110101100111", -- 15718 FREE #<CONS 0 15719>
 "00000000000000000011110101101000", -- 15719 FREE #<CONS 0 15720>
 "00000000000000000011110101101001", -- 15720 FREE #<CONS 0 15721>
 "00000000000000000011110101101010", -- 15721 FREE #<CONS 0 15722>
 "00000000000000000011110101101011", -- 15722 FREE #<CONS 0 15723>
 "00000000000000000011110101101100", -- 15723 FREE #<CONS 0 15724>
 "00000000000000000011110101101101", -- 15724 FREE #<CONS 0 15725>
 "00000000000000000011110101101110", -- 15725 FREE #<CONS 0 15726>
 "00000000000000000011110101101111", -- 15726 FREE #<CONS 0 15727>
 "00000000000000000011110101110000", -- 15727 FREE #<CONS 0 15728>
 "00000000000000000011110101110001", -- 15728 FREE #<CONS 0 15729>
 "00000000000000000011110101110010", -- 15729 FREE #<CONS 0 15730>
 "00000000000000000011110101110011", -- 15730 FREE #<CONS 0 15731>
 "00000000000000000011110101110100", -- 15731 FREE #<CONS 0 15732>
 "00000000000000000011110101110101", -- 15732 FREE #<CONS 0 15733>
 "00000000000000000011110101110110", -- 15733 FREE #<CONS 0 15734>
 "00000000000000000011110101110111", -- 15734 FREE #<CONS 0 15735>
 "00000000000000000011110101111000", -- 15735 FREE #<CONS 0 15736>
 "00000000000000000011110101111001", -- 15736 FREE #<CONS 0 15737>
 "00000000000000000011110101111010", -- 15737 FREE #<CONS 0 15738>
 "00000000000000000011110101111011", -- 15738 FREE #<CONS 0 15739>
 "00000000000000000011110101111100", -- 15739 FREE #<CONS 0 15740>
 "00000000000000000011110101111101", -- 15740 FREE #<CONS 0 15741>
 "00000000000000000011110101111110", -- 15741 FREE #<CONS 0 15742>
 "00000000000000000011110101111111", -- 15742 FREE #<CONS 0 15743>
 "00000000000000000011110110000000", -- 15743 FREE #<CONS 0 15744>
 "00000000000000000011110110000001", -- 15744 FREE #<CONS 0 15745>
 "00000000000000000011110110000010", -- 15745 FREE #<CONS 0 15746>
 "00000000000000000011110110000011", -- 15746 FREE #<CONS 0 15747>
 "00000000000000000011110110000100", -- 15747 FREE #<CONS 0 15748>
 "00000000000000000011110110000101", -- 15748 FREE #<CONS 0 15749>
 "00000000000000000011110110000110", -- 15749 FREE #<CONS 0 15750>
 "00000000000000000011110110000111", -- 15750 FREE #<CONS 0 15751>
 "00000000000000000011110110001000", -- 15751 FREE #<CONS 0 15752>
 "00000000000000000011110110001001", -- 15752 FREE #<CONS 0 15753>
 "00000000000000000011110110001010", -- 15753 FREE #<CONS 0 15754>
 "00000000000000000011110110001011", -- 15754 FREE #<CONS 0 15755>
 "00000000000000000011110110001100", -- 15755 FREE #<CONS 0 15756>
 "00000000000000000011110110001101", -- 15756 FREE #<CONS 0 15757>
 "00000000000000000011110110001110", -- 15757 FREE #<CONS 0 15758>
 "00000000000000000011110110001111", -- 15758 FREE #<CONS 0 15759>
 "00000000000000000011110110010000", -- 15759 FREE #<CONS 0 15760>
 "00000000000000000011110110010001", -- 15760 FREE #<CONS 0 15761>
 "00000000000000000011110110010010", -- 15761 FREE #<CONS 0 15762>
 "00000000000000000011110110010011", -- 15762 FREE #<CONS 0 15763>
 "00000000000000000011110110010100", -- 15763 FREE #<CONS 0 15764>
 "00000000000000000011110110010101", -- 15764 FREE #<CONS 0 15765>
 "00000000000000000011110110010110", -- 15765 FREE #<CONS 0 15766>
 "00000000000000000011110110010111", -- 15766 FREE #<CONS 0 15767>
 "00000000000000000011110110011000", -- 15767 FREE #<CONS 0 15768>
 "00000000000000000011110110011001", -- 15768 FREE #<CONS 0 15769>
 "00000000000000000011110110011010", -- 15769 FREE #<CONS 0 15770>
 "00000000000000000011110110011011", -- 15770 FREE #<CONS 0 15771>
 "00000000000000000011110110011100", -- 15771 FREE #<CONS 0 15772>
 "00000000000000000011110110011101", -- 15772 FREE #<CONS 0 15773>
 "00000000000000000011110110011110", -- 15773 FREE #<CONS 0 15774>
 "00000000000000000011110110011111", -- 15774 FREE #<CONS 0 15775>
 "00000000000000000011110110100000", -- 15775 FREE #<CONS 0 15776>
 "00000000000000000011110110100001", -- 15776 FREE #<CONS 0 15777>
 "00000000000000000011110110100010", -- 15777 FREE #<CONS 0 15778>
 "00000000000000000011110110100011", -- 15778 FREE #<CONS 0 15779>
 "00000000000000000011110110100100", -- 15779 FREE #<CONS 0 15780>
 "00000000000000000011110110100101", -- 15780 FREE #<CONS 0 15781>
 "00000000000000000011110110100110", -- 15781 FREE #<CONS 0 15782>
 "00000000000000000011110110100111", -- 15782 FREE #<CONS 0 15783>
 "00000000000000000011110110101000", -- 15783 FREE #<CONS 0 15784>
 "00000000000000000011110110101001", -- 15784 FREE #<CONS 0 15785>
 "00000000000000000011110110101010", -- 15785 FREE #<CONS 0 15786>
 "00000000000000000011110110101011", -- 15786 FREE #<CONS 0 15787>
 "00000000000000000011110110101100", -- 15787 FREE #<CONS 0 15788>
 "00000000000000000011110110101101", -- 15788 FREE #<CONS 0 15789>
 "00000000000000000011110110101110", -- 15789 FREE #<CONS 0 15790>
 "00000000000000000011110110101111", -- 15790 FREE #<CONS 0 15791>
 "00000000000000000011110110110000", -- 15791 FREE #<CONS 0 15792>
 "00000000000000000011110110110001", -- 15792 FREE #<CONS 0 15793>
 "00000000000000000011110110110010", -- 15793 FREE #<CONS 0 15794>
 "00000000000000000011110110110011", -- 15794 FREE #<CONS 0 15795>
 "00000000000000000011110110110100", -- 15795 FREE #<CONS 0 15796>
 "00000000000000000011110110110101", -- 15796 FREE #<CONS 0 15797>
 "00000000000000000011110110110110", -- 15797 FREE #<CONS 0 15798>
 "00000000000000000011110110110111", -- 15798 FREE #<CONS 0 15799>
 "00000000000000000011110110111000", -- 15799 FREE #<CONS 0 15800>
 "00000000000000000011110110111001", -- 15800 FREE #<CONS 0 15801>
 "00000000000000000011110110111010", -- 15801 FREE #<CONS 0 15802>
 "00000000000000000011110110111011", -- 15802 FREE #<CONS 0 15803>
 "00000000000000000011110110111100", -- 15803 FREE #<CONS 0 15804>
 "00000000000000000011110110111101", -- 15804 FREE #<CONS 0 15805>
 "00000000000000000011110110111110", -- 15805 FREE #<CONS 0 15806>
 "00000000000000000011110110111111", -- 15806 FREE #<CONS 0 15807>
 "00000000000000000011110111000000", -- 15807 FREE #<CONS 0 15808>
 "00000000000000000011110111000001", -- 15808 FREE #<CONS 0 15809>
 "00000000000000000011110111000010", -- 15809 FREE #<CONS 0 15810>
 "00000000000000000011110111000011", -- 15810 FREE #<CONS 0 15811>
 "00000000000000000011110111000100", -- 15811 FREE #<CONS 0 15812>
 "00000000000000000011110111000101", -- 15812 FREE #<CONS 0 15813>
 "00000000000000000011110111000110", -- 15813 FREE #<CONS 0 15814>
 "00000000000000000011110111000111", -- 15814 FREE #<CONS 0 15815>
 "00000000000000000011110111001000", -- 15815 FREE #<CONS 0 15816>
 "00000000000000000011110111001001", -- 15816 FREE #<CONS 0 15817>
 "00000000000000000011110111001010", -- 15817 FREE #<CONS 0 15818>
 "00000000000000000011110111001011", -- 15818 FREE #<CONS 0 15819>
 "00000000000000000011110111001100", -- 15819 FREE #<CONS 0 15820>
 "00000000000000000011110111001101", -- 15820 FREE #<CONS 0 15821>
 "00000000000000000011110111001110", -- 15821 FREE #<CONS 0 15822>
 "00000000000000000011110111001111", -- 15822 FREE #<CONS 0 15823>
 "00000000000000000011110111010000", -- 15823 FREE #<CONS 0 15824>
 "00000000000000000011110111010001", -- 15824 FREE #<CONS 0 15825>
 "00000000000000000011110111010010", -- 15825 FREE #<CONS 0 15826>
 "00000000000000000011110111010011", -- 15826 FREE #<CONS 0 15827>
 "00000000000000000011110111010100", -- 15827 FREE #<CONS 0 15828>
 "00000000000000000011110111010101", -- 15828 FREE #<CONS 0 15829>
 "00000000000000000011110111010110", -- 15829 FREE #<CONS 0 15830>
 "00000000000000000011110111010111", -- 15830 FREE #<CONS 0 15831>
 "00000000000000000011110111011000", -- 15831 FREE #<CONS 0 15832>
 "00000000000000000011110111011001", -- 15832 FREE #<CONS 0 15833>
 "00000000000000000011110111011010", -- 15833 FREE #<CONS 0 15834>
 "00000000000000000011110111011011", -- 15834 FREE #<CONS 0 15835>
 "00000000000000000011110111011100", -- 15835 FREE #<CONS 0 15836>
 "00000000000000000011110111011101", -- 15836 FREE #<CONS 0 15837>
 "00000000000000000011110111011110", -- 15837 FREE #<CONS 0 15838>
 "00000000000000000011110111011111", -- 15838 FREE #<CONS 0 15839>
 "00000000000000000011110111100000", -- 15839 FREE #<CONS 0 15840>
 "00000000000000000011110111100001", -- 15840 FREE #<CONS 0 15841>
 "00000000000000000011110111100010", -- 15841 FREE #<CONS 0 15842>
 "00000000000000000011110111100011", -- 15842 FREE #<CONS 0 15843>
 "00000000000000000011110111100100", -- 15843 FREE #<CONS 0 15844>
 "00000000000000000011110111100101", -- 15844 FREE #<CONS 0 15845>
 "00000000000000000011110111100110", -- 15845 FREE #<CONS 0 15846>
 "00000000000000000011110111100111", -- 15846 FREE #<CONS 0 15847>
 "00000000000000000011110111101000", -- 15847 FREE #<CONS 0 15848>
 "00000000000000000011110111101001", -- 15848 FREE #<CONS 0 15849>
 "00000000000000000011110111101010", -- 15849 FREE #<CONS 0 15850>
 "00000000000000000011110111101011", -- 15850 FREE #<CONS 0 15851>
 "00000000000000000011110111101100", -- 15851 FREE #<CONS 0 15852>
 "00000000000000000011110111101101", -- 15852 FREE #<CONS 0 15853>
 "00000000000000000011110111101110", -- 15853 FREE #<CONS 0 15854>
 "00000000000000000011110111101111", -- 15854 FREE #<CONS 0 15855>
 "00000000000000000011110111110000", -- 15855 FREE #<CONS 0 15856>
 "00000000000000000011110111110001", -- 15856 FREE #<CONS 0 15857>
 "00000000000000000011110111110010", -- 15857 FREE #<CONS 0 15858>
 "00000000000000000011110111110011", -- 15858 FREE #<CONS 0 15859>
 "00000000000000000011110111110100", -- 15859 FREE #<CONS 0 15860>
 "00000000000000000011110111110101", -- 15860 FREE #<CONS 0 15861>
 "00000000000000000011110111110110", -- 15861 FREE #<CONS 0 15862>
 "00000000000000000011110111110111", -- 15862 FREE #<CONS 0 15863>
 "00000000000000000011110111111000", -- 15863 FREE #<CONS 0 15864>
 "00000000000000000011110111111001", -- 15864 FREE #<CONS 0 15865>
 "00000000000000000011110111111010", -- 15865 FREE #<CONS 0 15866>
 "00000000000000000011110111111011", -- 15866 FREE #<CONS 0 15867>
 "00000000000000000011110111111100", -- 15867 FREE #<CONS 0 15868>
 "00000000000000000011110111111101", -- 15868 FREE #<CONS 0 15869>
 "00000000000000000011110111111110", -- 15869 FREE #<CONS 0 15870>
 "00000000000000000011110111111111", -- 15870 FREE #<CONS 0 15871>
 "00000000000000000011111000000000", -- 15871 FREE #<CONS 0 15872>
 "00000000000000000011111000000001", -- 15872 FREE #<CONS 0 15873>
 "00000000000000000011111000000010", -- 15873 FREE #<CONS 0 15874>
 "00000000000000000011111000000011", -- 15874 FREE #<CONS 0 15875>
 "00000000000000000011111000000100", -- 15875 FREE #<CONS 0 15876>
 "00000000000000000011111000000101", -- 15876 FREE #<CONS 0 15877>
 "00000000000000000011111000000110", -- 15877 FREE #<CONS 0 15878>
 "00000000000000000011111000000111", -- 15878 FREE #<CONS 0 15879>
 "00000000000000000011111000001000", -- 15879 FREE #<CONS 0 15880>
 "00000000000000000011111000001001", -- 15880 FREE #<CONS 0 15881>
 "00000000000000000011111000001010", -- 15881 FREE #<CONS 0 15882>
 "00000000000000000011111000001011", -- 15882 FREE #<CONS 0 15883>
 "00000000000000000011111000001100", -- 15883 FREE #<CONS 0 15884>
 "00000000000000000011111000001101", -- 15884 FREE #<CONS 0 15885>
 "00000000000000000011111000001110", -- 15885 FREE #<CONS 0 15886>
 "00000000000000000011111000001111", -- 15886 FREE #<CONS 0 15887>
 "00000000000000000011111000010000", -- 15887 FREE #<CONS 0 15888>
 "00000000000000000011111000010001", -- 15888 FREE #<CONS 0 15889>
 "00000000000000000011111000010010", -- 15889 FREE #<CONS 0 15890>
 "00000000000000000011111000010011", -- 15890 FREE #<CONS 0 15891>
 "00000000000000000011111000010100", -- 15891 FREE #<CONS 0 15892>
 "00000000000000000011111000010101", -- 15892 FREE #<CONS 0 15893>
 "00000000000000000011111000010110", -- 15893 FREE #<CONS 0 15894>
 "00000000000000000011111000010111", -- 15894 FREE #<CONS 0 15895>
 "00000000000000000011111000011000", -- 15895 FREE #<CONS 0 15896>
 "00000000000000000011111000011001", -- 15896 FREE #<CONS 0 15897>
 "00000000000000000011111000011010", -- 15897 FREE #<CONS 0 15898>
 "00000000000000000011111000011011", -- 15898 FREE #<CONS 0 15899>
 "00000000000000000011111000011100", -- 15899 FREE #<CONS 0 15900>
 "00000000000000000011111000011101", -- 15900 FREE #<CONS 0 15901>
 "00000000000000000011111000011110", -- 15901 FREE #<CONS 0 15902>
 "00000000000000000011111000011111", -- 15902 FREE #<CONS 0 15903>
 "00000000000000000011111000100000", -- 15903 FREE #<CONS 0 15904>
 "00000000000000000011111000100001", -- 15904 FREE #<CONS 0 15905>
 "00000000000000000011111000100010", -- 15905 FREE #<CONS 0 15906>
 "00000000000000000011111000100011", -- 15906 FREE #<CONS 0 15907>
 "00000000000000000011111000100100", -- 15907 FREE #<CONS 0 15908>
 "00000000000000000011111000100101", -- 15908 FREE #<CONS 0 15909>
 "00000000000000000011111000100110", -- 15909 FREE #<CONS 0 15910>
 "00000000000000000011111000100111", -- 15910 FREE #<CONS 0 15911>
 "00000000000000000011111000101000", -- 15911 FREE #<CONS 0 15912>
 "00000000000000000011111000101001", -- 15912 FREE #<CONS 0 15913>
 "00000000000000000011111000101010", -- 15913 FREE #<CONS 0 15914>
 "00000000000000000011111000101011", -- 15914 FREE #<CONS 0 15915>
 "00000000000000000011111000101100", -- 15915 FREE #<CONS 0 15916>
 "00000000000000000011111000101101", -- 15916 FREE #<CONS 0 15917>
 "00000000000000000011111000101110", -- 15917 FREE #<CONS 0 15918>
 "00000000000000000011111000101111", -- 15918 FREE #<CONS 0 15919>
 "00000000000000000011111000110000", -- 15919 FREE #<CONS 0 15920>
 "00000000000000000011111000110001", -- 15920 FREE #<CONS 0 15921>
 "00000000000000000011111000110010", -- 15921 FREE #<CONS 0 15922>
 "00000000000000000011111000110011", -- 15922 FREE #<CONS 0 15923>
 "00000000000000000011111000110100", -- 15923 FREE #<CONS 0 15924>
 "00000000000000000011111000110101", -- 15924 FREE #<CONS 0 15925>
 "00000000000000000011111000110110", -- 15925 FREE #<CONS 0 15926>
 "00000000000000000011111000110111", -- 15926 FREE #<CONS 0 15927>
 "00000000000000000011111000111000", -- 15927 FREE #<CONS 0 15928>
 "00000000000000000011111000111001", -- 15928 FREE #<CONS 0 15929>
 "00000000000000000011111000111010", -- 15929 FREE #<CONS 0 15930>
 "00000000000000000011111000111011", -- 15930 FREE #<CONS 0 15931>
 "00000000000000000011111000111100", -- 15931 FREE #<CONS 0 15932>
 "00000000000000000011111000111101", -- 15932 FREE #<CONS 0 15933>
 "00000000000000000011111000111110", -- 15933 FREE #<CONS 0 15934>
 "00000000000000000011111000111111", -- 15934 FREE #<CONS 0 15935>
 "00000000000000000011111001000000", -- 15935 FREE #<CONS 0 15936>
 "00000000000000000011111001000001", -- 15936 FREE #<CONS 0 15937>
 "00000000000000000011111001000010", -- 15937 FREE #<CONS 0 15938>
 "00000000000000000011111001000011", -- 15938 FREE #<CONS 0 15939>
 "00000000000000000011111001000100", -- 15939 FREE #<CONS 0 15940>
 "00000000000000000011111001000101", -- 15940 FREE #<CONS 0 15941>
 "00000000000000000011111001000110", -- 15941 FREE #<CONS 0 15942>
 "00000000000000000011111001000111", -- 15942 FREE #<CONS 0 15943>
 "00000000000000000011111001001000", -- 15943 FREE #<CONS 0 15944>
 "00000000000000000011111001001001", -- 15944 FREE #<CONS 0 15945>
 "00000000000000000011111001001010", -- 15945 FREE #<CONS 0 15946>
 "00000000000000000011111001001011", -- 15946 FREE #<CONS 0 15947>
 "00000000000000000011111001001100", -- 15947 FREE #<CONS 0 15948>
 "00000000000000000011111001001101", -- 15948 FREE #<CONS 0 15949>
 "00000000000000000011111001001110", -- 15949 FREE #<CONS 0 15950>
 "00000000000000000011111001001111", -- 15950 FREE #<CONS 0 15951>
 "00000000000000000011111001010000", -- 15951 FREE #<CONS 0 15952>
 "00000000000000000011111001010001", -- 15952 FREE #<CONS 0 15953>
 "00000000000000000011111001010010", -- 15953 FREE #<CONS 0 15954>
 "00000000000000000011111001010011", -- 15954 FREE #<CONS 0 15955>
 "00000000000000000011111001010100", -- 15955 FREE #<CONS 0 15956>
 "00000000000000000011111001010101", -- 15956 FREE #<CONS 0 15957>
 "00000000000000000011111001010110", -- 15957 FREE #<CONS 0 15958>
 "00000000000000000011111001010111", -- 15958 FREE #<CONS 0 15959>
 "00000000000000000011111001011000", -- 15959 FREE #<CONS 0 15960>
 "00000000000000000011111001011001", -- 15960 FREE #<CONS 0 15961>
 "00000000000000000011111001011010", -- 15961 FREE #<CONS 0 15962>
 "00000000000000000011111001011011", -- 15962 FREE #<CONS 0 15963>
 "00000000000000000011111001011100", -- 15963 FREE #<CONS 0 15964>
 "00000000000000000011111001011101", -- 15964 FREE #<CONS 0 15965>
 "00000000000000000011111001011110", -- 15965 FREE #<CONS 0 15966>
 "00000000000000000011111001011111", -- 15966 FREE #<CONS 0 15967>
 "00000000000000000011111001100000", -- 15967 FREE #<CONS 0 15968>
 "00000000000000000011111001100001", -- 15968 FREE #<CONS 0 15969>
 "00000000000000000011111001100010", -- 15969 FREE #<CONS 0 15970>
 "00000000000000000011111001100011", -- 15970 FREE #<CONS 0 15971>
 "00000000000000000011111001100100", -- 15971 FREE #<CONS 0 15972>
 "00000000000000000011111001100101", -- 15972 FREE #<CONS 0 15973>
 "00000000000000000011111001100110", -- 15973 FREE #<CONS 0 15974>
 "00000000000000000011111001100111", -- 15974 FREE #<CONS 0 15975>
 "00000000000000000011111001101000", -- 15975 FREE #<CONS 0 15976>
 "00000000000000000011111001101001", -- 15976 FREE #<CONS 0 15977>
 "00000000000000000011111001101010", -- 15977 FREE #<CONS 0 15978>
 "00000000000000000011111001101011", -- 15978 FREE #<CONS 0 15979>
 "00000000000000000011111001101100", -- 15979 FREE #<CONS 0 15980>
 "00000000000000000011111001101101", -- 15980 FREE #<CONS 0 15981>
 "00000000000000000011111001101110", -- 15981 FREE #<CONS 0 15982>
 "00000000000000000011111001101111", -- 15982 FREE #<CONS 0 15983>
 "00000000000000000011111001110000", -- 15983 FREE #<CONS 0 15984>
 "00000000000000000011111001110001", -- 15984 FREE #<CONS 0 15985>
 "00000000000000000011111001110010", -- 15985 FREE #<CONS 0 15986>
 "00000000000000000011111001110011", -- 15986 FREE #<CONS 0 15987>
 "00000000000000000011111001110100", -- 15987 FREE #<CONS 0 15988>
 "00000000000000000011111001110101", -- 15988 FREE #<CONS 0 15989>
 "00000000000000000011111001110110", -- 15989 FREE #<CONS 0 15990>
 "00000000000000000011111001110111", -- 15990 FREE #<CONS 0 15991>
 "00000000000000000011111001111000", -- 15991 FREE #<CONS 0 15992>
 "00000000000000000011111001111001", -- 15992 FREE #<CONS 0 15993>
 "00000000000000000011111001111010", -- 15993 FREE #<CONS 0 15994>
 "00000000000000000011111001111011", -- 15994 FREE #<CONS 0 15995>
 "00000000000000000011111001111100", -- 15995 FREE #<CONS 0 15996>
 "00000000000000000011111001111101", -- 15996 FREE #<CONS 0 15997>
 "00000000000000000011111001111110", -- 15997 FREE #<CONS 0 15998>
 "00000000000000000011111001111111", -- 15998 FREE #<CONS 0 15999>
 "00000000000000000011111010000000", -- 15999 FREE #<CONS 0 16000>
 "00000000000000000011111010000001", -- 16000 FREE #<CONS 0 16001>
 "00000000000000000011111010000010", -- 16001 FREE #<CONS 0 16002>
 "00000000000000000011111010000011", -- 16002 FREE #<CONS 0 16003>
 "00000000000000000011111010000100", -- 16003 FREE #<CONS 0 16004>
 "00000000000000000011111010000101", -- 16004 FREE #<CONS 0 16005>
 "00000000000000000011111010000110", -- 16005 FREE #<CONS 0 16006>
 "00000000000000000011111010000111", -- 16006 FREE #<CONS 0 16007>
 "00000000000000000011111010001000", -- 16007 FREE #<CONS 0 16008>
 "00000000000000000011111010001001", -- 16008 FREE #<CONS 0 16009>
 "00000000000000000011111010001010", -- 16009 FREE #<CONS 0 16010>
 "00000000000000000011111010001011", -- 16010 FREE #<CONS 0 16011>
 "00000000000000000011111010001100", -- 16011 FREE #<CONS 0 16012>
 "00000000000000000011111010001101", -- 16012 FREE #<CONS 0 16013>
 "00000000000000000011111010001110", -- 16013 FREE #<CONS 0 16014>
 "00000000000000000011111010001111", -- 16014 FREE #<CONS 0 16015>
 "00000000000000000011111010010000", -- 16015 FREE #<CONS 0 16016>
 "00000000000000000011111010010001", -- 16016 FREE #<CONS 0 16017>
 "00000000000000000011111010010010", -- 16017 FREE #<CONS 0 16018>
 "00000000000000000011111010010011", -- 16018 FREE #<CONS 0 16019>
 "00000000000000000011111010010100", -- 16019 FREE #<CONS 0 16020>
 "00000000000000000011111010010101", -- 16020 FREE #<CONS 0 16021>
 "00000000000000000011111010010110", -- 16021 FREE #<CONS 0 16022>
 "00000000000000000011111010010111", -- 16022 FREE #<CONS 0 16023>
 "00000000000000000011111010011000", -- 16023 FREE #<CONS 0 16024>
 "00000000000000000011111010011001", -- 16024 FREE #<CONS 0 16025>
 "00000000000000000011111010011010", -- 16025 FREE #<CONS 0 16026>
 "00000000000000000011111010011011", -- 16026 FREE #<CONS 0 16027>
 "00000000000000000011111010011100", -- 16027 FREE #<CONS 0 16028>
 "00000000000000000011111010011101", -- 16028 FREE #<CONS 0 16029>
 "00000000000000000011111010011110", -- 16029 FREE #<CONS 0 16030>
 "00000000000000000011111010011111", -- 16030 FREE #<CONS 0 16031>
 "00000000000000000011111010100000", -- 16031 FREE #<CONS 0 16032>
 "00000000000000000011111010100001", -- 16032 FREE #<CONS 0 16033>
 "00000000000000000011111010100010", -- 16033 FREE #<CONS 0 16034>
 "00000000000000000011111010100011", -- 16034 FREE #<CONS 0 16035>
 "00000000000000000011111010100100", -- 16035 FREE #<CONS 0 16036>
 "00000000000000000011111010100101", -- 16036 FREE #<CONS 0 16037>
 "00000000000000000011111010100110", -- 16037 FREE #<CONS 0 16038>
 "00000000000000000011111010100111", -- 16038 FREE #<CONS 0 16039>
 "00000000000000000011111010101000", -- 16039 FREE #<CONS 0 16040>
 "00000000000000000011111010101001", -- 16040 FREE #<CONS 0 16041>
 "00000000000000000011111010101010", -- 16041 FREE #<CONS 0 16042>
 "00000000000000000011111010101011", -- 16042 FREE #<CONS 0 16043>
 "00000000000000000011111010101100", -- 16043 FREE #<CONS 0 16044>
 "00000000000000000011111010101101", -- 16044 FREE #<CONS 0 16045>
 "00000000000000000011111010101110", -- 16045 FREE #<CONS 0 16046>
 "00000000000000000011111010101111", -- 16046 FREE #<CONS 0 16047>
 "00000000000000000011111010110000", -- 16047 FREE #<CONS 0 16048>
 "00000000000000000011111010110001", -- 16048 FREE #<CONS 0 16049>
 "00000000000000000011111010110010", -- 16049 FREE #<CONS 0 16050>
 "00000000000000000011111010110011", -- 16050 FREE #<CONS 0 16051>
 "00000000000000000011111010110100", -- 16051 FREE #<CONS 0 16052>
 "00000000000000000011111010110101", -- 16052 FREE #<CONS 0 16053>
 "00000000000000000011111010110110", -- 16053 FREE #<CONS 0 16054>
 "00000000000000000011111010110111", -- 16054 FREE #<CONS 0 16055>
 "00000000000000000011111010111000", -- 16055 FREE #<CONS 0 16056>
 "00000000000000000011111010111001", -- 16056 FREE #<CONS 0 16057>
 "00000000000000000011111010111010", -- 16057 FREE #<CONS 0 16058>
 "00000000000000000011111010111011", -- 16058 FREE #<CONS 0 16059>
 "00000000000000000011111010111100", -- 16059 FREE #<CONS 0 16060>
 "00000000000000000011111010111101", -- 16060 FREE #<CONS 0 16061>
 "00000000000000000011111010111110", -- 16061 FREE #<CONS 0 16062>
 "00000000000000000011111010111111", -- 16062 FREE #<CONS 0 16063>
 "00000000000000000011111011000000", -- 16063 FREE #<CONS 0 16064>
 "00000000000000000011111011000001", -- 16064 FREE #<CONS 0 16065>
 "00000000000000000011111011000010", -- 16065 FREE #<CONS 0 16066>
 "00000000000000000011111011000011", -- 16066 FREE #<CONS 0 16067>
 "00000000000000000011111011000100", -- 16067 FREE #<CONS 0 16068>
 "00000000000000000011111011000101", -- 16068 FREE #<CONS 0 16069>
 "00000000000000000011111011000110", -- 16069 FREE #<CONS 0 16070>
 "00000000000000000011111011000111", -- 16070 FREE #<CONS 0 16071>
 "00000000000000000011111011001000", -- 16071 FREE #<CONS 0 16072>
 "00000000000000000011111011001001", -- 16072 FREE #<CONS 0 16073>
 "00000000000000000011111011001010", -- 16073 FREE #<CONS 0 16074>
 "00000000000000000011111011001011", -- 16074 FREE #<CONS 0 16075>
 "00000000000000000011111011001100", -- 16075 FREE #<CONS 0 16076>
 "00000000000000000011111011001101", -- 16076 FREE #<CONS 0 16077>
 "00000000000000000011111011001110", -- 16077 FREE #<CONS 0 16078>
 "00000000000000000011111011001111", -- 16078 FREE #<CONS 0 16079>
 "00000000000000000011111011010000", -- 16079 FREE #<CONS 0 16080>
 "00000000000000000011111011010001", -- 16080 FREE #<CONS 0 16081>
 "00000000000000000011111011010010", -- 16081 FREE #<CONS 0 16082>
 "00000000000000000011111011010011", -- 16082 FREE #<CONS 0 16083>
 "00000000000000000011111011010100", -- 16083 FREE #<CONS 0 16084>
 "00000000000000000011111011010101", -- 16084 FREE #<CONS 0 16085>
 "00000000000000000011111011010110", -- 16085 FREE #<CONS 0 16086>
 "00000000000000000011111011010111", -- 16086 FREE #<CONS 0 16087>
 "00000000000000000011111011011000", -- 16087 FREE #<CONS 0 16088>
 "00000000000000000011111011011001", -- 16088 FREE #<CONS 0 16089>
 "00000000000000000011111011011010", -- 16089 FREE #<CONS 0 16090>
 "00000000000000000011111011011011", -- 16090 FREE #<CONS 0 16091>
 "00000000000000000011111011011100", -- 16091 FREE #<CONS 0 16092>
 "00000000000000000011111011011101", -- 16092 FREE #<CONS 0 16093>
 "00000000000000000011111011011110", -- 16093 FREE #<CONS 0 16094>
 "00000000000000000011111011011111", -- 16094 FREE #<CONS 0 16095>
 "00000000000000000011111011100000", -- 16095 FREE #<CONS 0 16096>
 "00000000000000000011111011100001", -- 16096 FREE #<CONS 0 16097>
 "00000000000000000011111011100010", -- 16097 FREE #<CONS 0 16098>
 "00000000000000000011111011100011", -- 16098 FREE #<CONS 0 16099>
 "00000000000000000011111011100100", -- 16099 FREE #<CONS 0 16100>
 "00000000000000000011111011100101", -- 16100 FREE #<CONS 0 16101>
 "00000000000000000011111011100110", -- 16101 FREE #<CONS 0 16102>
 "00000000000000000011111011100111", -- 16102 FREE #<CONS 0 16103>
 "00000000000000000011111011101000", -- 16103 FREE #<CONS 0 16104>
 "00000000000000000011111011101001", -- 16104 FREE #<CONS 0 16105>
 "00000000000000000011111011101010", -- 16105 FREE #<CONS 0 16106>
 "00000000000000000011111011101011", -- 16106 FREE #<CONS 0 16107>
 "00000000000000000011111011101100", -- 16107 FREE #<CONS 0 16108>
 "00000000000000000011111011101101", -- 16108 FREE #<CONS 0 16109>
 "00000000000000000011111011101110", -- 16109 FREE #<CONS 0 16110>
 "00000000000000000011111011101111", -- 16110 FREE #<CONS 0 16111>
 "00000000000000000011111011110000", -- 16111 FREE #<CONS 0 16112>
 "00000000000000000011111011110001", -- 16112 FREE #<CONS 0 16113>
 "00000000000000000011111011110010", -- 16113 FREE #<CONS 0 16114>
 "00000000000000000011111011110011", -- 16114 FREE #<CONS 0 16115>
 "00000000000000000011111011110100", -- 16115 FREE #<CONS 0 16116>
 "00000000000000000011111011110101", -- 16116 FREE #<CONS 0 16117>
 "00000000000000000011111011110110", -- 16117 FREE #<CONS 0 16118>
 "00000000000000000011111011110111", -- 16118 FREE #<CONS 0 16119>
 "00000000000000000011111011111000", -- 16119 FREE #<CONS 0 16120>
 "00000000000000000011111011111001", -- 16120 FREE #<CONS 0 16121>
 "00000000000000000011111011111010", -- 16121 FREE #<CONS 0 16122>
 "00000000000000000011111011111011", -- 16122 FREE #<CONS 0 16123>
 "00000000000000000011111011111100", -- 16123 FREE #<CONS 0 16124>
 "00000000000000000011111011111101", -- 16124 FREE #<CONS 0 16125>
 "00000000000000000011111011111110", -- 16125 FREE #<CONS 0 16126>
 "00000000000000000011111011111111", -- 16126 FREE #<CONS 0 16127>
 "00000000000000000011111100000000", -- 16127 FREE #<CONS 0 16128>
 "00000000000000000011111100000001", -- 16128 FREE #<CONS 0 16129>
 "00000000000000000011111100000010", -- 16129 FREE #<CONS 0 16130>
 "00000000000000000011111100000011", -- 16130 FREE #<CONS 0 16131>
 "00000000000000000011111100000100", -- 16131 FREE #<CONS 0 16132>
 "00000000000000000011111100000101", -- 16132 FREE #<CONS 0 16133>
 "00000000000000000011111100000110", -- 16133 FREE #<CONS 0 16134>
 "00000000000000000011111100000111", -- 16134 FREE #<CONS 0 16135>
 "00000000000000000011111100001000", -- 16135 FREE #<CONS 0 16136>
 "00000000000000000011111100001001", -- 16136 FREE #<CONS 0 16137>
 "00000000000000000011111100001010", -- 16137 FREE #<CONS 0 16138>
 "00000000000000000011111100001011", -- 16138 FREE #<CONS 0 16139>
 "00000000000000000011111100001100", -- 16139 FREE #<CONS 0 16140>
 "00000000000000000011111100001101", -- 16140 FREE #<CONS 0 16141>
 "00000000000000000011111100001110", -- 16141 FREE #<CONS 0 16142>
 "00000000000000000011111100001111", -- 16142 FREE #<CONS 0 16143>
 "00000000000000000011111100010000", -- 16143 FREE #<CONS 0 16144>
 "00000000000000000011111100010001", -- 16144 FREE #<CONS 0 16145>
 "00000000000000000011111100010010", -- 16145 FREE #<CONS 0 16146>
 "00000000000000000011111100010011", -- 16146 FREE #<CONS 0 16147>
 "00000000000000000011111100010100", -- 16147 FREE #<CONS 0 16148>
 "00000000000000000011111100010101", -- 16148 FREE #<CONS 0 16149>
 "00000000000000000011111100010110", -- 16149 FREE #<CONS 0 16150>
 "00000000000000000011111100010111", -- 16150 FREE #<CONS 0 16151>
 "00000000000000000011111100011000", -- 16151 FREE #<CONS 0 16152>
 "00000000000000000011111100011001", -- 16152 FREE #<CONS 0 16153>
 "00000000000000000011111100011010", -- 16153 FREE #<CONS 0 16154>
 "00000000000000000011111100011011", -- 16154 FREE #<CONS 0 16155>
 "00000000000000000011111100011100", -- 16155 FREE #<CONS 0 16156>
 "00000000000000000011111100011101", -- 16156 FREE #<CONS 0 16157>
 "00000000000000000011111100011110", -- 16157 FREE #<CONS 0 16158>
 "00000000000000000011111100011111", -- 16158 FREE #<CONS 0 16159>
 "00000000000000000011111100100000", -- 16159 FREE #<CONS 0 16160>
 "00000000000000000011111100100001", -- 16160 FREE #<CONS 0 16161>
 "00000000000000000011111100100010", -- 16161 FREE #<CONS 0 16162>
 "00000000000000000011111100100011", -- 16162 FREE #<CONS 0 16163>
 "00000000000000000011111100100100", -- 16163 FREE #<CONS 0 16164>
 "00000000000000000011111100100101", -- 16164 FREE #<CONS 0 16165>
 "00000000000000000011111100100110", -- 16165 FREE #<CONS 0 16166>
 "00000000000000000011111100100111", -- 16166 FREE #<CONS 0 16167>
 "00000000000000000011111100101000", -- 16167 FREE #<CONS 0 16168>
 "00000000000000000011111100101001", -- 16168 FREE #<CONS 0 16169>
 "00000000000000000011111100101010", -- 16169 FREE #<CONS 0 16170>
 "00000000000000000011111100101011", -- 16170 FREE #<CONS 0 16171>
 "00000000000000000011111100101100", -- 16171 FREE #<CONS 0 16172>
 "00000000000000000011111100101101", -- 16172 FREE #<CONS 0 16173>
 "00000000000000000011111100101110", -- 16173 FREE #<CONS 0 16174>
 "00000000000000000011111100101111", -- 16174 FREE #<CONS 0 16175>
 "00000000000000000011111100110000", -- 16175 FREE #<CONS 0 16176>
 "00000000000000000011111100110001", -- 16176 FREE #<CONS 0 16177>
 "00000000000000000011111100110010", -- 16177 FREE #<CONS 0 16178>
 "00000000000000000011111100110011", -- 16178 FREE #<CONS 0 16179>
 "00000000000000000011111100110100", -- 16179 FREE #<CONS 0 16180>
 "00000000000000000011111100110101", -- 16180 FREE #<CONS 0 16181>
 "00000000000000000011111100110110", -- 16181 FREE #<CONS 0 16182>
 "00000000000000000011111100110111", -- 16182 FREE #<CONS 0 16183>
 "00000000000000000011111100111000", -- 16183 FREE #<CONS 0 16184>
 "00000000000000000011111100111001", -- 16184 FREE #<CONS 0 16185>
 "00000000000000000011111100111010", -- 16185 FREE #<CONS 0 16186>
 "00000000000000000011111100111011", -- 16186 FREE #<CONS 0 16187>
 "00000000000000000011111100111100", -- 16187 FREE #<CONS 0 16188>
 "00000000000000000011111100111101", -- 16188 FREE #<CONS 0 16189>
 "00000000000000000011111100111110", -- 16189 FREE #<CONS 0 16190>
 "00000000000000000011111100111111", -- 16190 FREE #<CONS 0 16191>
 "00000000000000000011111101000000", -- 16191 FREE #<CONS 0 16192>
 "00000000000000000011111101000001", -- 16192 FREE #<CONS 0 16193>
 "00000000000000000011111101000010", -- 16193 FREE #<CONS 0 16194>
 "00000000000000000011111101000011", -- 16194 FREE #<CONS 0 16195>
 "00000000000000000011111101000100", -- 16195 FREE #<CONS 0 16196>
 "00000000000000000011111101000101", -- 16196 FREE #<CONS 0 16197>
 "00000000000000000011111101000110", -- 16197 FREE #<CONS 0 16198>
 "00000000000000000011111101000111", -- 16198 FREE #<CONS 0 16199>
 "00000000000000000011111101001000", -- 16199 FREE #<CONS 0 16200>
 "00000000000000000011111101001001", -- 16200 FREE #<CONS 0 16201>
 "00000000000000000011111101001010", -- 16201 FREE #<CONS 0 16202>
 "00000000000000000011111101001011", -- 16202 FREE #<CONS 0 16203>
 "00000000000000000011111101001100", -- 16203 FREE #<CONS 0 16204>
 "00000000000000000011111101001101", -- 16204 FREE #<CONS 0 16205>
 "00000000000000000011111101001110", -- 16205 FREE #<CONS 0 16206>
 "00000000000000000011111101001111", -- 16206 FREE #<CONS 0 16207>
 "00000000000000000011111101010000", -- 16207 FREE #<CONS 0 16208>
 "00000000000000000011111101010001", -- 16208 FREE #<CONS 0 16209>
 "00000000000000000011111101010010", -- 16209 FREE #<CONS 0 16210>
 "00000000000000000011111101010011", -- 16210 FREE #<CONS 0 16211>
 "00000000000000000011111101010100", -- 16211 FREE #<CONS 0 16212>
 "00000000000000000011111101010101", -- 16212 FREE #<CONS 0 16213>
 "00000000000000000011111101010110", -- 16213 FREE #<CONS 0 16214>
 "00000000000000000011111101010111", -- 16214 FREE #<CONS 0 16215>
 "00000000000000000011111101011000", -- 16215 FREE #<CONS 0 16216>
 "00000000000000000011111101011001", -- 16216 FREE #<CONS 0 16217>
 "00000000000000000011111101011010", -- 16217 FREE #<CONS 0 16218>
 "00000000000000000011111101011011", -- 16218 FREE #<CONS 0 16219>
 "00000000000000000011111101011100", -- 16219 FREE #<CONS 0 16220>
 "00000000000000000011111101011101", -- 16220 FREE #<CONS 0 16221>
 "00000000000000000011111101011110", -- 16221 FREE #<CONS 0 16222>
 "00000000000000000011111101011111", -- 16222 FREE #<CONS 0 16223>
 "00000000000000000011111101100000", -- 16223 FREE #<CONS 0 16224>
 "00000000000000000011111101100001", -- 16224 FREE #<CONS 0 16225>
 "00000000000000000011111101100010", -- 16225 FREE #<CONS 0 16226>
 "00000000000000000011111101100011", -- 16226 FREE #<CONS 0 16227>
 "00000000000000000011111101100100", -- 16227 FREE #<CONS 0 16228>
 "00000000000000000011111101100101", -- 16228 FREE #<CONS 0 16229>
 "00000000000000000011111101100110", -- 16229 FREE #<CONS 0 16230>
 "00000000000000000011111101100111", -- 16230 FREE #<CONS 0 16231>
 "00000000000000000011111101101000", -- 16231 FREE #<CONS 0 16232>
 "00000000000000000011111101101001", -- 16232 FREE #<CONS 0 16233>
 "00000000000000000011111101101010", -- 16233 FREE #<CONS 0 16234>
 "00000000000000000011111101101011", -- 16234 FREE #<CONS 0 16235>
 "00000000000000000011111101101100", -- 16235 FREE #<CONS 0 16236>
 "00000000000000000011111101101101", -- 16236 FREE #<CONS 0 16237>
 "00000000000000000011111101101110", -- 16237 FREE #<CONS 0 16238>
 "00000000000000000011111101101111", -- 16238 FREE #<CONS 0 16239>
 "00000000000000000011111101110000", -- 16239 FREE #<CONS 0 16240>
 "00000000000000000011111101110001", -- 16240 FREE #<CONS 0 16241>
 "00000000000000000011111101110010", -- 16241 FREE #<CONS 0 16242>
 "00000000000000000011111101110011", -- 16242 FREE #<CONS 0 16243>
 "00000000000000000011111101110100", -- 16243 FREE #<CONS 0 16244>
 "00000000000000000011111101110101", -- 16244 FREE #<CONS 0 16245>
 "00000000000000000011111101110110", -- 16245 FREE #<CONS 0 16246>
 "00000000000000000011111101110111", -- 16246 FREE #<CONS 0 16247>
 "00000000000000000011111101111000", -- 16247 FREE #<CONS 0 16248>
 "00000000000000000011111101111001", -- 16248 FREE #<CONS 0 16249>
 "00000000000000000011111101111010", -- 16249 FREE #<CONS 0 16250>
 "00000000000000000011111101111011", -- 16250 FREE #<CONS 0 16251>
 "00000000000000000011111101111100", -- 16251 FREE #<CONS 0 16252>
 "00000000000000000011111101111101", -- 16252 FREE #<CONS 0 16253>
 "00000000000000000011111101111110", -- 16253 FREE #<CONS 0 16254>
 "00000000000000000011111101111111", -- 16254 FREE #<CONS 0 16255>
 "00000000000000000011111110000000", -- 16255 FREE #<CONS 0 16256>
 "00000000000000000011111110000001", -- 16256 FREE #<CONS 0 16257>
 "00000000000000000011111110000010", -- 16257 FREE #<CONS 0 16258>
 "00000000000000000011111110000011", -- 16258 FREE #<CONS 0 16259>
 "00000000000000000011111110000100", -- 16259 FREE #<CONS 0 16260>
 "00000000000000000011111110000101", -- 16260 FREE #<CONS 0 16261>
 "00000000000000000011111110000110", -- 16261 FREE #<CONS 0 16262>
 "00000000000000000011111110000111", -- 16262 FREE #<CONS 0 16263>
 "00000000000000000011111110001000", -- 16263 FREE #<CONS 0 16264>
 "00000000000000000011111110001001", -- 16264 FREE #<CONS 0 16265>
 "00000000000000000011111110001010", -- 16265 FREE #<CONS 0 16266>
 "00000000000000000011111110001011", -- 16266 FREE #<CONS 0 16267>
 "00000000000000000011111110001100", -- 16267 FREE #<CONS 0 16268>
 "00000000000000000011111110001101", -- 16268 FREE #<CONS 0 16269>
 "00000000000000000011111110001110", -- 16269 FREE #<CONS 0 16270>
 "00000000000000000011111110001111", -- 16270 FREE #<CONS 0 16271>
 "00000000000000000011111110010000", -- 16271 FREE #<CONS 0 16272>
 "00000000000000000011111110010001", -- 16272 FREE #<CONS 0 16273>
 "00000000000000000011111110010010", -- 16273 FREE #<CONS 0 16274>
 "00000000000000000011111110010011", -- 16274 FREE #<CONS 0 16275>
 "00000000000000000011111110010100", -- 16275 FREE #<CONS 0 16276>
 "00000000000000000011111110010101", -- 16276 FREE #<CONS 0 16277>
 "00000000000000000011111110010110", -- 16277 FREE #<CONS 0 16278>
 "00000000000000000011111110010111", -- 16278 FREE #<CONS 0 16279>
 "00000000000000000011111110011000", -- 16279 FREE #<CONS 0 16280>
 "00000000000000000011111110011001", -- 16280 FREE #<CONS 0 16281>
 "00000000000000000011111110011010", -- 16281 FREE #<CONS 0 16282>
 "00000000000000000011111110011011", -- 16282 FREE #<CONS 0 16283>
 "00000000000000000011111110011100", -- 16283 FREE #<CONS 0 16284>
 "00000000000000000011111110011101", -- 16284 FREE #<CONS 0 16285>
 "00000000000000000011111110011110", -- 16285 FREE #<CONS 0 16286>
 "00000000000000000011111110011111", -- 16286 FREE #<CONS 0 16287>
 "00000000000000000011111110100000", -- 16287 FREE #<CONS 0 16288>
 "00000000000000000011111110100001", -- 16288 FREE #<CONS 0 16289>
 "00000000000000000011111110100010", -- 16289 FREE #<CONS 0 16290>
 "00000000000000000011111110100011", -- 16290 FREE #<CONS 0 16291>
 "00000000000000000011111110100100", -- 16291 FREE #<CONS 0 16292>
 "00000000000000000011111110100101", -- 16292 FREE #<CONS 0 16293>
 "00000000000000000011111110100110", -- 16293 FREE #<CONS 0 16294>
 "00000000000000000011111110100111", -- 16294 FREE #<CONS 0 16295>
 "00000000000000000011111110101000", -- 16295 FREE #<CONS 0 16296>
 "00000000000000000011111110101001", -- 16296 FREE #<CONS 0 16297>
 "00000000000000000011111110101010", -- 16297 FREE #<CONS 0 16298>
 "00000000000000000011111110101011", -- 16298 FREE #<CONS 0 16299>
 "00000000000000000011111110101100", -- 16299 FREE #<CONS 0 16300>
 "00000000000000000011111110101101", -- 16300 FREE #<CONS 0 16301>
 "00000000000000000011111110101110", -- 16301 FREE #<CONS 0 16302>
 "00000000000000000011111110101111", -- 16302 FREE #<CONS 0 16303>
 "00000000000000000011111110110000", -- 16303 FREE #<CONS 0 16304>
 "00000000000000000011111110110001", -- 16304 FREE #<CONS 0 16305>
 "00000000000000000011111110110010", -- 16305 FREE #<CONS 0 16306>
 "00000000000000000011111110110011", -- 16306 FREE #<CONS 0 16307>
 "00000000000000000011111110110100", -- 16307 FREE #<CONS 0 16308>
 "00000000000000000011111110110101", -- 16308 FREE #<CONS 0 16309>
 "00000000000000000011111110110110", -- 16309 FREE #<CONS 0 16310>
 "00000000000000000011111110110111", -- 16310 FREE #<CONS 0 16311>
 "00000000000000000011111110111000", -- 16311 FREE #<CONS 0 16312>
 "00000000000000000011111110111001", -- 16312 FREE #<CONS 0 16313>
 "00000000000000000011111110111010", -- 16313 FREE #<CONS 0 16314>
 "00000000000000000011111110111011", -- 16314 FREE #<CONS 0 16315>
 "00000000000000000011111110111100", -- 16315 FREE #<CONS 0 16316>
 "00000000000000000011111110111101", -- 16316 FREE #<CONS 0 16317>
 "00000000000000000011111110111110", -- 16317 FREE #<CONS 0 16318>
 "00000000000000000011111110111111", -- 16318 FREE #<CONS 0 16319>
 "00000000000000000011111111000000", -- 16319 FREE #<CONS 0 16320>
 "00000000000000000011111111000001", -- 16320 FREE #<CONS 0 16321>
 "00000000000000000011111111000010", -- 16321 FREE #<CONS 0 16322>
 "00000000000000000011111111000011", -- 16322 FREE #<CONS 0 16323>
 "00000000000000000011111111000100", -- 16323 FREE #<CONS 0 16324>
 "00000000000000000011111111000101", -- 16324 FREE #<CONS 0 16325>
 "00000000000000000011111111000110", -- 16325 FREE #<CONS 0 16326>
 "00000000000000000011111111000111", -- 16326 FREE #<CONS 0 16327>
 "00000000000000000011111111001000", -- 16327 FREE #<CONS 0 16328>
 "00000000000000000011111111001001", -- 16328 FREE #<CONS 0 16329>
 "00000000000000000011111111001010", -- 16329 FREE #<CONS 0 16330>
 "00000000000000000011111111001011", -- 16330 FREE #<CONS 0 16331>
 "00000000000000000011111111001100", -- 16331 FREE #<CONS 0 16332>
 "00000000000000000011111111001101", -- 16332 FREE #<CONS 0 16333>
 "00000000000000000011111111001110", -- 16333 FREE #<CONS 0 16334>
 "00000000000000000011111111001111", -- 16334 FREE #<CONS 0 16335>
 "00000000000000000011111111010000", -- 16335 FREE #<CONS 0 16336>
 "00000000000000000011111111010001", -- 16336 FREE #<CONS 0 16337>
 "00000000000000000011111111010010", -- 16337 FREE #<CONS 0 16338>
 "00000000000000000011111111010011", -- 16338 FREE #<CONS 0 16339>
 "00000000000000000011111111010100", -- 16339 FREE #<CONS 0 16340>
 "00000000000000000011111111010101", -- 16340 FREE #<CONS 0 16341>
 "00000000000000000011111111010110", -- 16341 FREE #<CONS 0 16342>
 "00000000000000000011111111010111", -- 16342 FREE #<CONS 0 16343>
 "00000000000000000011111111011000", -- 16343 FREE #<CONS 0 16344>
 "00000000000000000011111111011001", -- 16344 FREE #<CONS 0 16345>
 "00000000000000000011111111011010", -- 16345 FREE #<CONS 0 16346>
 "00000000000000000011111111011011", -- 16346 FREE #<CONS 0 16347>
 "00000000000000000011111111011100", -- 16347 FREE #<CONS 0 16348>
 "00000000000000000011111111011101", -- 16348 FREE #<CONS 0 16349>
 "00000000000000000011111111011110", -- 16349 FREE #<CONS 0 16350>
 "00000000000000000011111111011111", -- 16350 FREE #<CONS 0 16351>
 "00000000000000000011111111100000", -- 16351 FREE #<CONS 0 16352>
 "00000000000000000011111111100001", -- 16352 FREE #<CONS 0 16353>
 "00000000000000000011111111100010", -- 16353 FREE #<CONS 0 16354>
 "00000000000000000011111111100011", -- 16354 FREE #<CONS 0 16355>
 "00000000000000000011111111100100", -- 16355 FREE #<CONS 0 16356>
 "00000000000000000011111111100101", -- 16356 FREE #<CONS 0 16357>
 "00000000000000000011111111100110", -- 16357 FREE #<CONS 0 16358>
 "00000000000000000011111111100111", -- 16358 FREE #<CONS 0 16359>
 "00000000000000000011111111101000", -- 16359 FREE #<CONS 0 16360>
 "00000000000000000011111111101001", -- 16360 FREE #<CONS 0 16361>
 "00000000000000000011111111101010", -- 16361 FREE #<CONS 0 16362>
 "00000000000000000011111111101011", -- 16362 FREE #<CONS 0 16363>
 "00000000000000000011111111101100", -- 16363 FREE #<CONS 0 16364>
 "00000000000000000011111111101101", -- 16364 FREE #<CONS 0 16365>
 "00000000000000000011111111101110", -- 16365 FREE #<CONS 0 16366>
 "00000000000000000011111111101111", -- 16366 FREE #<CONS 0 16367>
 "00000000000000000011111111110000", -- 16367 FREE #<CONS 0 16368>
 "00000000000000000011111111110001", -- 16368 FREE #<CONS 0 16369>
 "00000000000000000011111111110010", -- 16369 FREE #<CONS 0 16370>
 "00000000000000000011111111110011", -- 16370 FREE #<CONS 0 16371>
 "00000000000000000011111111110100", -- 16371 FREE #<CONS 0 16372>
 "00000000000000000011111111110101", -- 16372 FREE #<CONS 0 16373>
 "00000000000000000011111111110110", -- 16373 FREE #<CONS 0 16374>
 "00000000000000000011111111110111", -- 16374 FREE #<CONS 0 16375>
 "00000000000000000011111111111000", -- 16375 FREE #<CONS 0 16376>
 "00000000000000000011111111111001", -- 16376 FREE #<CONS 0 16377>
 "00000000000000000011111111111010", -- 16377 FREE #<CONS 0 16378>
 "00000000000000000011111111111011", -- 16378 FREE #<CONS 0 16379>
 "00000000000000000011111111111100", -- 16379 FREE #<CONS 0 16380>
 "00000000000000000011111111111101", -- 16380 FREE #<CONS 0 16381>
 "00000000000000000011111111111110", -- 16381 FREE #<CONS 0 16382>
 "00000000000000000011111111111111", -- 16382 FREE #<CONS 0 16383>
 "00000000101110011000001011100111" -- 16383 INITIALIZE #<CONS 742 743>
);

end package;

