--
-- KBUG9S
-- 4 September 2004
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
library unisim;
use unisim.all;

entity mon_rom is
  Port (
    clk   : in  std_logic;
    cs    : in  std_logic;
    addr  : in  std_logic_vector (10 downto 0);
    rdata : out std_logic_vector (7 downto 0)
    );
end mon_rom;

architecture rtl of mon_rom is

  component RAMB16_S9
    generic (
      INIT_00, INIT_01, INIT_02, INIT_03,
      INIT_04, INIT_05, INIT_06, INIT_07,
      INIT_08, INIT_09, INIT_0A, INIT_0B,
      INIT_0C, INIT_0D, INIT_0E, INIT_0F,
      INIT_10, INIT_11, INIT_12, INIT_13,
      INIT_14, INIT_15, INIT_16, INIT_17,
      INIT_18, INIT_19, INIT_1A, INIT_1B,
      INIT_1C, INIT_1D, INIT_1E, INIT_1F,
      INIT_20, INIT_21, INIT_22, INIT_23,
      INIT_24, INIT_25, INIT_26, INIT_27,
      INIT_28, INIT_29, INIT_2A, INIT_2B,
      INIT_2C, INIT_2D, INIT_2E, INIT_2F,
      INIT_30, INIT_31, INIT_32, INIT_33,
      INIT_34, INIT_35, INIT_36, INIT_37,
      INIT_38, INIT_39, INIT_3A, INIT_3B,
      INIT_3C, INIT_3D, INIT_3E, INIT_3F : bit_vector (255 downto 0)
      );

    port (
      do   : out std_logic_vector(7 downto 0);
      dop  : out std_logic_vector(0 downto 0);
      addr : in std_logic_vector(10 downto 0);
      clk  : in std_logic;
      di   : in std_logic_vector(7 downto 0);
      dip  : in std_logic_vector(0 downto 0);
      we   : in std_logic;
      en   : in std_logic;
      ssr  : in std_logic
      );
  end component RAMB16_S9;

  signal dp : std_logic;

begin

  ROM : RAMB16_S9
    generic map (
      INIT_00 => x"FBFC1BFD18FA18FA18FA18FA18FA4FFC53FC5EFCABFC65FCA9FC80FC7CF838F8",
      INIT_01 => x"C6C0F08E10B9FE8EC0F0CE100CFD04FDFBFCFAFCEBFCDCFCD2FCBFFC3AFD04FD",
      INIT_02 => x"A7D0866AAFDD8C30FB265AE26F0CC68E0117D0F0BF00E08EF9265AA0A780A610",
      -- INIT_03 => x"17E5FE8EE20317C9FE8EA504178704174F0417D8F0B70A86D7F0B70386431FE4", -- (unpatched)
      INIT_03 => x"1700007EE20317C9FE8EA504178704174F0417D8F0B70A86D7F0B70386431FE4", -- (patched)
      INIT_04 => x"A302170E0417408B981F1504175E86092C2081891FF1270D817F84FB0317CD03",
      INIT_05 => x"1F2D29450217C22094ADC620AA0317E7FE8EF526B9FE8C02300F2780E17AFE8E",
      INIT_06 => x"E127088111283802176C0217650317A4A6740217650317211F880317EDFE8E12",
      INIT_07 => x"31C2202131B003173F864D02170827A4A1A4A7390F260D8117275E81DD271881",
      INIT_08 => x"1000C3101F390124E1AC20340629E6011705201F30C0F08E321FC00217BE203F",
      INIT_09 => x"E4AE110317EDFE8E103439623203273403170527E4AC011FF0C4201F0634F0C4",
      INIT_0a => x"0425208180A610C6E1AEEB0117F5265AF30117EC021780A610C6FB0117EE0217",
      INIT_0b => x"17072653810503175F3B341F390128FD0117BC20EE265A4203172E8602237E81",
      INIT_0c => x"1F031707265381E702175F39D7F0F7E72001C88E031707265681F22002D83D03",
      INIT_0d => x"8E10341A24C0F08C1E294C011739D8F0F7E72008C84F031707264B81F22002D8",
      INIT_0e => x"10CC02163F866901173984A73F86A4AFA0A709273F8184A60F271035558DFFFF",
      INIT_0f => x"AE7DFE16AC0117068D4AAF0427268D1F304AAE431F39FB265A188D08C6D9F08E",
      INIT_10 => x"A608C6D9F08E1039A0A7A0A7A0A7FF8684A7A4A604263F8184A60A24C0F08C21",
      INIT_11 => x"273981670217F92653816E0217D2F07F528D1186393D3139F7265A0427A1ACA0",
      INIT_12 => x"170434E46AE46AE4EBE0EBE0E610342129B3001726290234CA0017F12631813C",
      INIT_13 => x"D2F073058D3F86B327FFC102355FEB2080A70527E46AE0EB02340C290435B000",
      INIT_14 => x"062762A3E4EC1102171286E4AF0130462562AC4A2930346F8DE26F2602161386",
      INIT_15 => x"63EB62EB75011762AE820117981F03CB9F01172EFF8E64E720C6022320008310",
      INIT_16 => x"188D3965326A8D1486C326E4AC62AF680117981F53F526646A72011780A684EB",
      INIT_17 => x"2D86121F4229088D391035F726E4AC1080A7A0A60929188D5D8D3E8610341529",
      INIT_18 => x"1E29078D891F484848482829118D903561A710343229088D011F38290E8D438D",
      INIT_19 => x"021A393780032246810725418139308003223981122530817C011739E0AB0434",
      INIT_1a => x"3941A70229B78DEA8D8300173944AF0229B38DF68D8500176301162086008D39",
      INIT_1b => x"AF0229858DC88D7C8D394AAF0229908DD38D7E8D3943A70229AB8DDE8D800017",
      INIT_1c => x"FF17A58D748D3942A702297DFF17B18D778D3946AF022979FF17BD8D7A8D3948",
      INIT_1d => x"358D910017EDFE8E348D2D8D268D1E8D168DA10017EDFE8E39C4A7808A042971",
      INIT_1e => x"A67F8D15FF8E572044AE88001709FF8E6120311F920017F1FE8E4A20438D3C8D",
      INIT_1f => x"FF8E332048AE648DFDFE8E3C204AAE6D8DF7FE8E4D2043A6768D0FFF8E562041",
      INIT_20 => x"80A608C6023426FF8EC4A6498D1FFF8E292042A6528D1AFF8E2A2046AE5B8D03",
      INIT_21 => x"8D4444444402340235028D023510348235EF265A17FF178200172D860225E468",
      INIT_22 => x"80A64D8D9035048DDFFE8E10340B20028D5C20078B022F3981308B0F84023504",
      INIT_23 => x"86354F0126800017052708C54F0B26618D042702C54FD8F0F6063439F8260481",
      INIT_24 => x"022066001705276200170A2708C510204C00170527478D092702C5D8F0F60434",
      INIT_25 => x"BE84357D0017032701C5358D022702C5D7F0F60434D58DD727D2F07D8435E020",
      INIT_26 => x"F0BE103482350185D0F09FA6023439D2F0B7FF86016D84A7118684A70386D0F0",
      INIT_27 => x"10E0B6023439943501A7FA2702C584E6D0F0BE1434903501A6FA27018584A6D0",
      INIT_28 => x"00CC20E08E943501A7FA2702C584E610E08E14343911E0B6FC27F58D82350185",
      INIT_29 => x"7D20E08E16345986028D1B86D6F07F01E702C6D5F0FD04E703E702A7D3F0FD00",
      INIT_2a => x"101B814100271008819635C5001784A70520098D042420810D20748D0427D6F0",
      INIT_2b => x"0027100B812C0027100C81990027100D814500271016818E0027101A816C0027",
      INIT_2c => x"F0B67400165A3C0027105DD3F0FC9900168300261019C15CD3F0FC51260A8111",
      INIT_2d => x"273DC1D6F0F65800160000CC5B00162500271050814CD3F0B66800164A3327D3",
      INIT_2e => x"39D5F0B70426D5F07D39D6F07F39D6F0B704263D81312754816E002710598116",
      INIT_2f => x"C6D3F0B6168D0000CC1B20E12218C120C0D5F07FD5F0F6ED224F812080D6F07F",
      INIT_30 => x"50814CD3F0FC3903E702A7D3F0FDD4F0F64F39D6F07FF726508102A74C84E720",
      INIT_31 => x"A702E7D3F0F72086D3F0F604E75F012519C15C04E6E78D5AEA2619C15C4FF026",
      INIT_32 => x"39D6F0F702E7D3F0F75FE4205F03E7D4F0F7082719C15CD4F0F6F42650C15C84",
      INIT_33 => x"8EFB0254FB01E62073FE178FFE17EE20CAFE176FFE17F6276AFE170D2698FE17",
      INIT_34 => x"F9496EF9470FF945B3F94260FE4182FB1948FB1877FB156CFB1060FB049AFB03",
      INIT_35 => x"F976F976F976F9DEFA5ADFF95803F953A8FB5285FA5077F94FBAF84D2CFA4C95",
      INIT_36 => x"0D0420302E31562053394755422D4B0000000A0D000000FFFFFFFFEBF976F976",
      INIT_37 => x"552020043D43502020043D5053202004202D20043F54414857043E040000000A",
      INIT_38 => x"20043D422020043D412020043D50442020043D58492020043D59492020043D50",
      INIT_39 => x"00000000000000000000000000000004315343565A4E4948464504203A434320",
      INIT_3a => x"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3b => x"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3c => x"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3d => x"9F6EC6F09F6EC4F09F6EC0F09F6E000000000000000000000000000000000000",
      INIT_3e => x"0822CEF0BC8B300F27FFFF8CCCF0BE49584F4AAF80E64AAE431FCAF09F6EC8F0",
      INIT_3f => x"34F834F8C2FFBEFFBAFFB6FFC6FFB2FFC2F09F6E42EE1F37F16E44AEC4EC1034"
      )

    port map (
      do   => rdata,
      dop(0) => dp,
      addr => addr,
      clk  => clk,
      dip(0) => dp,
      ssr => '0',
      di => (others => '0'),
      en   => cs,
      we   => '0'
      );

end architecture rtl;

